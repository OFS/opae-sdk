// ed_sim.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module ed_sim (
		output wire         ddr4a_waitrequest_n, //         ddr4a.waitrequest_n
		input  wire         ddr4a_read,          //              .read
		input  wire         ddr4a_write,         //              .write
		input  wire [25:0]  ddr4a_address,       //              .address
		output wire [511:0] ddr4a_readdata,      //              .readdata
		input  wire [511:0] ddr4a_writedata,     //              .writedata
		input  wire [6:0]   ddr4a_burstcount,    //              .burstcount
		input  wire [63:0]  ddr4a_byteenable,    //              .byteenable
		output wire         ddr4a_readdatavalid, //              .readdatavalid
		output wire         ddr4a_userclk_clk,   // ddr4a_userclk.clk
		output wire         ddr4b_waitrequest_n, //         ddr4b.waitrequest_n
		input  wire         ddr4b_read,          //              .read
		input  wire         ddr4b_write,         //              .write
		input  wire [25:0]  ddr4b_address,       //              .address
		output wire [511:0] ddr4b_readdata,      //              .readdata
		input  wire [511:0] ddr4b_writedata,     //              .writedata
		input  wire [6:0]   ddr4b_burstcount,    //              .burstcount
		input  wire [63:0]  ddr4b_byteenable,    //              .byteenable
		output wire         ddr4b_readdatavalid  //              .readdatavalid
	);

	wire         ed_sim_clock_source_0_clk_clk;                      // ed_sim_clock_source_0:clk -> [ddr4a:pll_ref_clk, ed_sim_reset_source_0:clk]
	wire  [31:0] ddr4a_clks_sharing_master_out_clks_sharing;         // ddr4a:clks_sharing_master_out -> clks_sharing_splitter:sig_input
	wire   [0:0] ddr4a_mem_mem_reset_n;                              // ddr4a:mem_reset_n -> mem_a:mem_reset_n
	wire   [1:0] ddr4a_mem_mem_ba;                                   // ddr4a:mem_ba -> mem_a:mem_ba
	wire   [1:0] ddr4a_mem_mem_bg;                                   // ddr4a:mem_bg -> mem_a:mem_bg
	wire   [0:0] ddr4a_mem_mem_ck;                                   // ddr4a:mem_ck -> mem_a:mem_ck
	wire   [7:0] ddr4a_mem_mem_dqs;                                  // [] -> [ddr4a:mem_dqs, mem_a:mem_dqs]
	wire   [0:0] ddr4a_mem_mem_act_n;                                // ddr4a:mem_act_n -> mem_a:mem_act_n
	wire  [63:0] ddr4a_mem_mem_dq;                                   // [] -> [ddr4a:mem_dq, mem_a:mem_dq]
	wire   [0:0] ddr4a_mem_mem_cs_n;                                 // ddr4a:mem_cs_n -> mem_a:mem_cs_n
	wire  [16:0] ddr4a_mem_mem_a;                                    // ddr4a:mem_a -> mem_a:mem_a
	wire   [0:0] ddr4a_mem_mem_odt;                                  // ddr4a:mem_odt -> mem_a:mem_odt
	wire   [0:0] mem_a_mem_mem_alert_n;                              // mem_a:mem_alert_n -> ddr4a:mem_alert_n
	wire   [7:0] ddr4a_mem_mem_dqs_n;                                // [] -> [ddr4a:mem_dqs_n, mem_a:mem_dqs_n]
	wire   [0:0] ddr4a_mem_mem_par;                                  // ddr4a:mem_par -> mem_a:mem_par
	wire   [7:0] ddr4a_mem_mem_dbi_n;                                // [] -> [ddr4a:mem_dbi_n, mem_a:mem_dbi_n]
	wire   [0:0] ddr4a_mem_mem_ck_n;                                 // ddr4a:mem_ck_n -> mem_a:mem_ck_n
	wire   [0:0] ddr4a_mem_mem_cke;                                  // ddr4a:mem_cke -> mem_a:mem_cke
	wire   [0:0] ddr4b_mem_mem_reset_n;                              // ddr4b:mem_reset_n -> mem_b:mem_reset_n
	wire   [1:0] ddr4b_mem_mem_ba;                                   // ddr4b:mem_ba -> mem_b:mem_ba
	wire   [1:0] ddr4b_mem_mem_bg;                                   // ddr4b:mem_bg -> mem_b:mem_bg
	wire   [0:0] ddr4b_mem_mem_ck;                                   // ddr4b:mem_ck -> mem_b:mem_ck
	wire   [7:0] ddr4b_mem_mem_dqs;                                  // [] -> [ddr4b:mem_dqs, mem_b:mem_dqs]
	wire   [0:0] ddr4b_mem_mem_act_n;                                // ddr4b:mem_act_n -> mem_b:mem_act_n
	wire  [63:0] ddr4b_mem_mem_dq;                                   // [] -> [ddr4b:mem_dq, mem_b:mem_dq]
	wire   [0:0] ddr4b_mem_mem_cs_n;                                 // ddr4b:mem_cs_n -> mem_b:mem_cs_n
	wire  [16:0] ddr4b_mem_mem_a;                                    // ddr4b:mem_a -> mem_b:mem_a
	wire   [0:0] ddr4b_mem_mem_odt;                                  // ddr4b:mem_odt -> mem_b:mem_odt
	wire   [0:0] mem_b_mem_mem_alert_n;                              // mem_b:mem_alert_n -> ddr4b:mem_alert_n
	wire   [7:0] ddr4b_mem_mem_dqs_n;                                // [] -> [ddr4b:mem_dqs_n, mem_b:mem_dqs_n]
	wire   [0:0] ddr4b_mem_mem_par;                                  // ddr4b:mem_par -> mem_b:mem_par
	wire   [7:0] ddr4b_mem_mem_dbi_n;                                // [] -> [ddr4b:mem_dbi_n, mem_b:mem_dbi_n]
	wire   [0:0] ddr4b_mem_mem_ck_n;                                 // ddr4b:mem_ck_n -> mem_b:mem_ck_n
	wire   [0:0] ddr4b_mem_mem_cke;                                  // ddr4b:mem_cke -> mem_b:mem_cke
	wire  [31:0] clks_sharing_splitter_sig_output_if_0_clks_sharing; // clks_sharing_splitter:sig_output_0 -> ddr4b:clks_sharing_slave_in
	wire         ed_sim_reset_source_0_reset_reset;                  // ed_sim_reset_source_0:reset -> ddr4a:global_reset_n

	ed_sim_clks_sharing_splitter clks_sharing_splitter (
		.sig_input    (ddr4a_clks_sharing_master_out_clks_sharing),         //    sig_input_if.clks_sharing
		.sig_output_0 (clks_sharing_splitter_sig_output_if_0_clks_sharing)  // sig_output_if_0.clks_sharing
	);

	ed_sim_ddr4a ddr4a (
		.clks_sharing_master_out (ddr4a_clks_sharing_master_out_clks_sharing), // clks_sharing_master_out.clks_sharing
		.amm_ready_0             (ddr4a_waitrequest_n),                        //              ctrl_amm_0.waitrequest_n
		.amm_read_0              (ddr4a_read),                                 //                        .read
		.amm_write_0             (ddr4a_write),                                //                        .write
		.amm_address_0           (ddr4a_address),                              //                        .address
		.amm_readdata_0          (ddr4a_readdata),                             //                        .readdata
		.amm_writedata_0         (ddr4a_writedata),                            //                        .writedata
		.amm_burstcount_0        (ddr4a_burstcount),                           //                        .burstcount
		.amm_byteenable_0        (ddr4a_byteenable),                           //                        .byteenable
		.amm_readdatavalid_0     (ddr4a_readdatavalid),                        //                        .readdatavalid
		.emif_usr_clk            (ddr4a_userclk_clk),                          //            emif_usr_clk.clk
		.emif_usr_reset_n        (),                                           //        emif_usr_reset_n.reset_n
		.global_reset_n          (ed_sim_reset_source_0_reset_reset),          //          global_reset_n.reset_n
		.mem_ck                  (ddr4a_mem_mem_ck),                           //                     mem.mem_ck
		.mem_ck_n                (ddr4a_mem_mem_ck_n),                         //                        .mem_ck_n
		.mem_a                   (ddr4a_mem_mem_a),                            //                        .mem_a
		.mem_act_n               (ddr4a_mem_mem_act_n),                        //                        .mem_act_n
		.mem_ba                  (ddr4a_mem_mem_ba),                           //                        .mem_ba
		.mem_bg                  (ddr4a_mem_mem_bg),                           //                        .mem_bg
		.mem_cke                 (ddr4a_mem_mem_cke),                          //                        .mem_cke
		.mem_cs_n                (ddr4a_mem_mem_cs_n),                         //                        .mem_cs_n
		.mem_odt                 (ddr4a_mem_mem_odt),                          //                        .mem_odt
		.mem_reset_n             (ddr4a_mem_mem_reset_n),                      //                        .mem_reset_n
		.mem_par                 (ddr4a_mem_mem_par),                          //                        .mem_par
		.mem_alert_n             (mem_a_mem_mem_alert_n),                      //                        .mem_alert_n
		.mem_dqs                 (ddr4a_mem_mem_dqs),                          //                        .mem_dqs
		.mem_dqs_n               (ddr4a_mem_mem_dqs_n),                        //                        .mem_dqs_n
		.mem_dq                  (ddr4a_mem_mem_dq),                           //                        .mem_dq
		.mem_dbi_n               (ddr4a_mem_mem_dbi_n),                        //                        .mem_dbi_n
		.oct_rzqin               (),                                           //                     oct.oct_rzqin
		.pll_ref_clk             (ed_sim_clock_source_0_clk_clk),              //             pll_ref_clk.clk
		.local_cal_success       (),                                           //                  status.local_cal_success
		.local_cal_fail          ()                                            //                        .local_cal_fail
	);

	ed_sim_emif_slave_1 ddr4b (
		.clks_sharing_slave_in (clks_sharing_splitter_sig_output_if_0_clks_sharing), // clks_sharing_slave_in.clks_sharing
		.amm_ready_0           (ddr4b_waitrequest_n),                                //            ctrl_amm_0.waitrequest_n
		.amm_read_0            (ddr4b_read),                                         //                      .read
		.amm_write_0           (ddr4b_write),                                        //                      .write
		.amm_address_0         (ddr4b_address),                                      //                      .address
		.amm_readdata_0        (ddr4b_readdata),                                     //                      .readdata
		.amm_writedata_0       (ddr4b_writedata),                                    //                      .writedata
		.amm_burstcount_0      (ddr4b_burstcount),                                   //                      .burstcount
		.amm_byteenable_0      (ddr4b_byteenable),                                   //                      .byteenable
		.amm_readdatavalid_0   (ddr4b_readdatavalid),                                //                      .readdatavalid
		.emif_usr_clk          (),                                                   //          emif_usr_clk.clk
		.emif_usr_reset_n      (),                                                   //      emif_usr_reset_n.reset_n
		.mem_ck                (ddr4b_mem_mem_ck),                                   //                   mem.mem_ck
		.mem_ck_n              (ddr4b_mem_mem_ck_n),                                 //                      .mem_ck_n
		.mem_a                 (ddr4b_mem_mem_a),                                    //                      .mem_a
		.mem_act_n             (ddr4b_mem_mem_act_n),                                //                      .mem_act_n
		.mem_ba                (ddr4b_mem_mem_ba),                                   //                      .mem_ba
		.mem_bg                (ddr4b_mem_mem_bg),                                   //                      .mem_bg
		.mem_cke               (ddr4b_mem_mem_cke),                                  //                      .mem_cke
		.mem_cs_n              (ddr4b_mem_mem_cs_n),                                 //                      .mem_cs_n
		.mem_odt               (ddr4b_mem_mem_odt),                                  //                      .mem_odt
		.mem_reset_n           (ddr4b_mem_mem_reset_n),                              //                      .mem_reset_n
		.mem_par               (ddr4b_mem_mem_par),                                  //                      .mem_par
		.mem_alert_n           (mem_b_mem_mem_alert_n),                              //                      .mem_alert_n
		.mem_dqs               (ddr4b_mem_mem_dqs),                                  //                      .mem_dqs
		.mem_dqs_n             (ddr4b_mem_mem_dqs_n),                                //                      .mem_dqs_n
		.mem_dq                (ddr4b_mem_mem_dq),                                   //                      .mem_dq
		.mem_dbi_n             (ddr4b_mem_mem_dbi_n),                                //                      .mem_dbi_n
		.oct_rzqin             (),                                                   //                   oct.oct_rzqin
		.local_cal_success     (),                                                   //                status.local_cal_success
		.local_cal_fail        ()                                                    //                      .local_cal_fail
	);

	ed_sim_pll_ref_clk_source ed_sim_clock_source_0 (
		.clk (ed_sim_clock_source_0_clk_clk)  // clk.clk
	);

	ed_sim_global_reset_n_source ed_sim_reset_source_0 (
		.clk   (ed_sim_clock_source_0_clk_clk),     //   clk.clk
		.reset (ed_sim_reset_source_0_reset_reset)  // reset.reset_n
	);

	ed_sim_mem_0 mem_a (
		.mem_ck      (ddr4a_mem_mem_ck),      // mem.mem_ck
		.mem_ck_n    (ddr4a_mem_mem_ck_n),    //    .mem_ck_n
		.mem_a       (ddr4a_mem_mem_a),       //    .mem_a
		.mem_act_n   (ddr4a_mem_mem_act_n),   //    .mem_act_n
		.mem_ba      (ddr4a_mem_mem_ba),      //    .mem_ba
		.mem_bg      (ddr4a_mem_mem_bg),      //    .mem_bg
		.mem_cke     (ddr4a_mem_mem_cke),     //    .mem_cke
		.mem_cs_n    (ddr4a_mem_mem_cs_n),    //    .mem_cs_n
		.mem_odt     (ddr4a_mem_mem_odt),     //    .mem_odt
		.mem_reset_n (ddr4a_mem_mem_reset_n), //    .mem_reset_n
		.mem_par     (ddr4a_mem_mem_par),     //    .mem_par
		.mem_alert_n (mem_a_mem_mem_alert_n), //    .mem_alert_n
		.mem_dqs     (ddr4a_mem_mem_dqs),     //    .mem_dqs
		.mem_dqs_n   (ddr4a_mem_mem_dqs_n),   //    .mem_dqs_n
		.mem_dq      (ddr4a_mem_mem_dq),      //    .mem_dq
		.mem_dbi_n   (ddr4a_mem_mem_dbi_n)    //    .mem_dbi_n
	);

	ed_sim_mem_1 mem_b (
		.mem_ck      (ddr4b_mem_mem_ck),      // mem.mem_ck
		.mem_ck_n    (ddr4b_mem_mem_ck_n),    //    .mem_ck_n
		.mem_a       (ddr4b_mem_mem_a),       //    .mem_a
		.mem_act_n   (ddr4b_mem_mem_act_n),   //    .mem_act_n
		.mem_ba      (ddr4b_mem_mem_ba),      //    .mem_ba
		.mem_bg      (ddr4b_mem_mem_bg),      //    .mem_bg
		.mem_cke     (ddr4b_mem_mem_cke),     //    .mem_cke
		.mem_cs_n    (ddr4b_mem_mem_cs_n),    //    .mem_cs_n
		.mem_odt     (ddr4b_mem_mem_odt),     //    .mem_odt
		.mem_reset_n (ddr4b_mem_mem_reset_n), //    .mem_reset_n
		.mem_par     (ddr4b_mem_mem_par),     //    .mem_par
		.mem_alert_n (mem_b_mem_mem_alert_n), //    .mem_alert_n
		.mem_dqs     (ddr4b_mem_mem_dqs),     //    .mem_dqs
		.mem_dqs_n   (ddr4b_mem_mem_dqs_n),   //    .mem_dqs_n
		.mem_dq      (ddr4b_mem_mem_dq),      //    .mem_dq
		.mem_dbi_n   (ddr4b_mem_mem_dbi_n)    //    .mem_dbi_n
	);

endmodule
