// ed_sim_global_reset_n_splitter.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module ed_sim_global_reset_n_splitter (
		input  wire  sig_input,    //    sig_input_if.reset_n
		output wire  sig_output_0  // sig_output_if_0.reset_n
	);

	assign sig_output_0 = sig_input;

endmodule
