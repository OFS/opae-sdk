// ed_sim_mem_0.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module ed_sim_mem_0 (
		input  wire [0:0]  mem_ck,      // mem.mem_ck
		input  wire [0:0]  mem_ck_n,    //    .mem_ck_n
		input  wire [16:0] mem_a,       //    .mem_a
		input  wire [0:0]  mem_act_n,   //    .mem_act_n
		input  wire [1:0]  mem_ba,      //    .mem_ba
		input  wire [1:0]  mem_bg,      //    .mem_bg
		input  wire [0:0]  mem_cke,     //    .mem_cke
		input  wire [0:0]  mem_cs_n,    //    .mem_cs_n
		input  wire [0:0]  mem_odt,     //    .mem_odt
		input  wire [0:0]  mem_reset_n, //    .mem_reset_n
		input  wire [0:0]  mem_par,     //    .mem_par
		output wire [0:0]  mem_alert_n, //    .mem_alert_n
		inout  wire [7:0]  mem_dqs,     //    .mem_dqs
		inout  wire [7:0]  mem_dqs_n,   //    .mem_dqs_n
		inout  wire [63:0] mem_dq,      //    .mem_dq
		inout  wire [7:0]  mem_dbi_n    //    .mem_dbi_n
	);

	ed_sim_mem_0_altera_emif_mem_model_170_nzcko3q mem_0 (
		.mem_ck      (mem_ck),      // mem.mem_ck
		.mem_ck_n    (mem_ck_n),    //    .mem_ck_n
		.mem_a       (mem_a),       //    .mem_a
		.mem_act_n   (mem_act_n),   //    .mem_act_n
		.mem_ba      (mem_ba),      //    .mem_ba
		.mem_bg      (mem_bg),      //    .mem_bg
		.mem_cke     (mem_cke),     //    .mem_cke
		.mem_cs_n    (mem_cs_n),    //    .mem_cs_n
		.mem_odt     (mem_odt),     //    .mem_odt
		.mem_reset_n (mem_reset_n), //    .mem_reset_n
		.mem_par     (mem_par),     //    .mem_par
		.mem_alert_n (mem_alert_n), //    .mem_alert_n
		.mem_dqs     (mem_dqs),     //    .mem_dqs
		.mem_dqs_n   (mem_dqs_n),   //    .mem_dqs_n
		.mem_dq      (mem_dq),      //    .mem_dq
		.mem_dbi_n   (mem_dbi_n)    //    .mem_dbi_n
	);

endmodule
