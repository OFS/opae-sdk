// ed_sim_global_reset_n_source.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module ed_sim_global_reset_n_source (
		input  wire  clk,   //   clk.clk
		output wire  reset  // reset.reset_n
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (5)
	) global_reset_n_source (
		.reset (reset), // reset.reset_n
		.clk   (clk)    //   clk.clk
	);

endmodule
