// (C) 2001-2017 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other
// Redistribution  and  use  in source  and  binary  forms,  with  or  without
// modification, are permitted provided that the following conditions are met:
//
// * Redistributions of  source code  must retain the  above copyright notice,
//   this list of conditions and the following disclaimer.
// * Redistributions in binary form must reproduce the above copyright notice,
//   this list of conditions and the following disclaimer in the documentation
//   and/or other materials provided with the distribution.
// * Neither the name  of Intel Corporation  nor the names of its contributors
//   may be used to  endorse or promote  products derived  from this  software
//   without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING,  BUT NOT LIMITED TO,  THE
// IMPLIED WARRANTIES OF  MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED.  IN NO EVENT  SHALL THE COPYRIGHT OWNER  OR CONTRIBUTORS BE
// LIABLE  FOR  ANY  DIRECT,  INDIRECT,  INCIDENTAL,  SPECIAL,  EXEMPLARY,  OR
// CONSEQUENTIAL  DAMAGES  (INCLUDING,  BUT  NOT LIMITED  TO,  PROCUREMENT  OF
// SUBSTITUTE GOODS OR SERVICES;  LOSS OF USE,  DATA, OR PROFITS;  OR BUSINESS
// INTERRUPTION)  HOWEVER CAUSED  AND ON ANY THEORY  OF LIABILITY,  WHETHER IN
// CONTRACT,  STRICT LIABILITY,  OR TORT  (INCLUDING NEGLIGENCE  OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE,  EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.



module io_12_lane_bcm__nf5es_abphy (
	ac_hmc,
	afi_rlat_core,
	afi_wlat_core,
	atbi_0,
	atbi_1,
	atpg_en_n,
	avl_address_in,
	avl_address_out,
	avl_clk_in,
	avl_clk_out,
	avl_read_in,
	avl_read_out,
	avl_readdata_in,
	avl_readdata_out,
	avl_write_in,
	avl_write_out,
	avl_writedata_in,
	avl_writedata_out,
	bhniotri,
	broadcast_in_bot,
	broadcast_in_top,
	broadcast_out_bot,
	broadcast_out_top,
	cas_csrdin,
	cas_csrdout,
	cfg_cmd_rate,
	cfg_dbc_ctrl_sel,
	cfg_dbc_dualport_en,
	cfg_dbc_in_protocol,
	cfg_dbc_pipe_lat,
	cfg_dbc_rc_en,
	cfg_dbc_slot_offset,
	cfg_dbc_slot_rotate_en,
	cfg_output_regd,
	cfg_reorder_rdata,
	cfg_rmw_en,
	clk_pll,
	codin_n,
	codin_nb,
	codin_p,
	codin_pb,
	core2dbc_rd_data_rdy,
	core2dbc_wr_data_vld0,
	core2dbc_wr_data_vld1,
	core2dbc_wr_ecc_info,
	core_dll,
	crnt_clk,
	csr_clk,
	csr_clk_left,
	csr_en,
	csr_en_left,
	csr_in,
	csr_out,
	csr_shift_n,
	ctl2dbc_cs0,
	ctl2dbc_cs1,
	ctl2dbc_mask_entry0,
	ctl2dbc_mask_entry1,
	ctl2dbc_misc0,
	ctl2dbc_misc1,
	ctl2dbc_mrnk_read0,
	ctl2dbc_mrnk_read1,
	ctl2dbc_nop0,
	ctl2dbc_nop1,
	ctl2dbc_rb_rdptr0,
	ctl2dbc_rb_rdptr1,
	ctl2dbc_rb_rdptr_vld0,
	ctl2dbc_rb_rdptr_vld1,
	ctl2dbc_rb_wrptr0,
	ctl2dbc_rb_wrptr1,
	ctl2dbc_rb_wrptr_vld0,
	ctl2dbc_rb_wrptr_vld1,
	ctl2dbc_rd_type0,
	ctl2dbc_rd_type1,
	ctl2dbc_rdata_en_full0,
	ctl2dbc_rdata_en_full1,
	ctl2dbc_seq_en0,
	ctl2dbc_seq_en1,
	ctl2dbc_wb_rdptr0,
	ctl2dbc_wb_rdptr1,
	ctl2dbc_wb_rdptr_vld0,
	ctl2dbc_wb_rdptr_vld1,
	ctl2dbc_wrdata_vld0,
	ctl2dbc_wrdata_vld1,
	data_from_core,
	data_to_core,
	dbc2core_rd_data_vld0,
	dbc2core_rd_data_vld1,
	dbc2core_rd_type,
	dbc2core_wb_pointer,
	dbc2core_wr_data_rdy,
	dbc2ctl_all_rd_done,
	dbc2ctl_rb_retire_ptr,
	dbc2ctl_rb_retire_ptr_vld,
	dbc2ctl_rd_data_vld,
	dbc2ctl_wb_retire_ptr,
	dbc2ctl_wb_retire_ptr_vld,
	dbc2db_wb_wrptr,
	dbc2db_wb_wrptr_vld,
	dft_core2db,
	dft_db2core,
	dft_phy_clk,
	dft_prbs_done,
	dft_prbs_ena_n,
	dft_prbs_pass,
	dll_core,
	dq_diff_in,
	dq_sstl_in,
	dqs_diff_in_0,
	dqs_diff_in_1,
	dqs_diff_in_2,
	dqs_diff_in_3,
	dqs_sstl_n_0,
	dqs_sstl_n_1,
	dqs_sstl_n_2,
	dqs_sstl_n_3,
	dqs_sstl_p_0,
	dqs_sstl_p_1,
	dqs_sstl_p_2,
	dqs_sstl_p_3,
	dzoutx,
	early_bhniotri,
	early_csren,
	early_enrnsl,
	early_frzreg,
	early_nfrzdrv,
	early_niotri,
	early_plniotri,
	early_usrmode,
	enrnsl,
	entest,
	fb_clkout,
	fr_in_clk,
	fr_out_clk,
	frzreg,
	hps_to_core_ctrl_en,
	hr_in_clk,
	hr_out_clk,
	i50u_ref,
	ibp50u,
	ibp50u_cal,
	ioereg_locked,
	jtag_clk,
	jtag_highz,
	jtag_mode,
	jtag_sdin,
	jtag_sdout,
	jtag_shftdr,
	jtag_updtdr,
	lane_cal_done,
	local_bhniotri,
	local_enrnsl,
	local_frzreg,
	local_nfrzdrv,
	local_niotri,
	local_plniotri,
	local_usrmode,
	local_wkpullup,
	lvds_rx_clk_chnl0,
	lvds_rx_clk_chnl1,
	lvds_rx_clk_chnl2,
	lvds_rx_clk_chnl3,
	lvds_rx_clk_chnl4,
	lvds_rx_clk_chnl5,
	lvds_tx_clk_chnl0,
	lvds_tx_clk_chnl1,
	lvds_tx_clk_chnl2,
	lvds_tx_clk_chnl3,
	lvds_tx_clk_chnl4,
	lvds_tx_clk_chnl5,
	mrnk_read_core,
	mrnk_write_core,
	n_crnt_clk,
	n_next_clk,
	naclr,
	ncein,
	nceout,
	next_clk,
	nfrzdrv,
	niotri,
	nsclr,
	oct_enable,
	oeb_from_core,
	osc_en_n,
	osc_enable_in,
	osc_mode_in,
	osc_rocount_to_core,
	osc_sel_n,
	phy_clk,
	phy_clk_phs,
	pipeline_global_en_n,
	pll_clk,
	pll_locked,
	plniotri,
	progctl,
	progoe,
	progout,
	rdata_en_full_core,
	rdata_valid_core,
	regulator_clk,
	reinit,
	reset_n,
	scan_shift_n,
	scanin,
	scanout,
	switch_dn,
	switch_up,
	sync_clk_bot_in,
	sync_clk_bot_out,
	sync_clk_top_in,
	sync_clk_top_out,
	sync_data_bot_in,
	sync_data_bot_out,
	sync_data_top_in,
	sync_data_top_out,
	test_avl_clk_in_en_n,
	test_clk,
	test_clk_ph_buf_en_n,
	test_clk_pll_en_n,
	test_clr_n,
	test_datovr_en_n,
	test_db_csr_in,
	test_dbg_in,
	test_dbg_out,
	test_dqs_csr_in,
	test_dqs_enable_en_n,
	test_fr_clk_en_n,
	test_hr_clk_en_n,
	test_int_clk_en_n,
	test_interp_clk_en_n,
	test_ioereg2_csr_out,
	test_phy_clk_en_n,
	test_phy_clk_lane_en_n,
	test_pst_clk_en_n,
	test_pst_dll_i,
	test_pst_dll_o,
	test_tdf_select_n,
	test_vref_csr_out,
	test_xor_clk,
	tpctl,
	tpdata,
	tpin,
	up_ph,
	usrmode,
	vref_ext,
	vref_int,
	weak_pullup_enable,
	wkpullup,
	x1024_osc_out,
	xor_vref,
	xprio_clk,
	xprio_sync,
	xprio_xbus
);

  timeunit 1ps;
  timeprecision 1ps;


	input [95:0]	ac_hmc;
	output [5:0]	afi_rlat_core;
	output [5:0]	afi_wlat_core;
	output	atbi_0;
	output	atbi_1;
	input	atpg_en_n;
	input [19:0]	avl_address_in;
	output [19:0]	avl_address_out;
	input	avl_clk_in;
	output	avl_clk_out;
	input	avl_read_in;
	output	avl_read_out;
	input [31:0]	avl_readdata_in;
	output [31:0]	avl_readdata_out;
	input	avl_write_in;
	output	avl_write_out;
	input [31:0]	avl_writedata_in;
	output [31:0]	avl_writedata_out;
	input	bhniotri;
	input	broadcast_in_bot;
	input	broadcast_in_top;
	output	broadcast_out_bot;
	output	broadcast_out_top;
	input [4:0]	cas_csrdin;
	output [4:0]	cas_csrdout;
	input [2:0]	cfg_cmd_rate;
	input	cfg_dbc_ctrl_sel;
	input	cfg_dbc_dualport_en;
	input	cfg_dbc_in_protocol;
	input [2:0]	cfg_dbc_pipe_lat;
	input	cfg_dbc_rc_en;
	input [1:0]	cfg_dbc_slot_offset;
	input [2:0]	cfg_dbc_slot_rotate_en;
	input	cfg_output_regd;
	input	cfg_reorder_rdata;
	input	cfg_rmw_en;
	input	clk_pll;
	output [11:0]	codin_n;
	output [11:0]	codin_nb;
	output [11:0]	codin_p;
	output [11:0]	codin_pb;
	input	core2dbc_rd_data_rdy;
	input	core2dbc_wr_data_vld0;
	input	core2dbc_wr_data_vld1;
	input [12:0]	core2dbc_wr_ecc_info;
	input [2:0]	core_dll;
	output [5:0]	crnt_clk;
	input	csr_clk;
	output	csr_clk_left;
	input	csr_en;
	output	csr_en_left;
	input	csr_in;
	output	csr_out;
	input	csr_shift_n;
	input [1:0]	ctl2dbc_cs0;
	input [1:0]	ctl2dbc_cs1;
	input	ctl2dbc_mask_entry0;
	input	ctl2dbc_mask_entry1;
	input [3:0]	ctl2dbc_misc0;
	input [3:0]	ctl2dbc_misc1;
	input [7:0]	ctl2dbc_mrnk_read0;
	input [7:0]	ctl2dbc_mrnk_read1;
	input	ctl2dbc_nop0;
	input	ctl2dbc_nop1;
	input [11:0]	ctl2dbc_rb_rdptr0;
	input [11:0]	ctl2dbc_rb_rdptr1;
	input [1:0]	ctl2dbc_rb_rdptr_vld0;
	input [1:0]	ctl2dbc_rb_rdptr_vld1;
	input [5:0]	ctl2dbc_rb_wrptr0;
	input [5:0]	ctl2dbc_rb_wrptr1;
	input	ctl2dbc_rb_wrptr_vld0;
	input	ctl2dbc_rb_wrptr_vld1;
	input	ctl2dbc_rd_type0;
	input	ctl2dbc_rd_type1;
	input [3:0]	ctl2dbc_rdata_en_full0;
	input [3:0]	ctl2dbc_rdata_en_full1;
	input	ctl2dbc_seq_en0;
	input	ctl2dbc_seq_en1;
	input [5:0]	ctl2dbc_wb_rdptr0;
	input [5:0]	ctl2dbc_wb_rdptr1;
	input	ctl2dbc_wb_rdptr_vld0;
	input	ctl2dbc_wb_rdptr_vld1;
	input	ctl2dbc_wrdata_vld0;
	input	ctl2dbc_wrdata_vld1;
	input [95:0]	data_from_core;
	output [95:0]	data_to_core;
	output	dbc2core_rd_data_vld0;
	output	dbc2core_rd_data_vld1;
	output	dbc2core_rd_type;
	output [11:0]	dbc2core_wb_pointer;
	output	dbc2core_wr_data_rdy;
	output	dbc2ctl_all_rd_done;
	output [5:0]	dbc2ctl_rb_retire_ptr;
	output	dbc2ctl_rb_retire_ptr_vld;
	output	dbc2ctl_rd_data_vld;
	output [5:0]	dbc2ctl_wb_retire_ptr;
	output	dbc2ctl_wb_retire_ptr_vld;
	output [5:0]	dbc2db_wb_wrptr;
	output	dbc2db_wb_wrptr_vld;
	input [7:0]	dft_core2db;
	output [7:0]	dft_db2core;
	output [1:0]	dft_phy_clk;
	output	dft_prbs_done;
	input	dft_prbs_ena_n;
	output	dft_prbs_pass;
	output [12:0]	dll_core;
	input [23:0]	dq_diff_in;
	input [23:0]	dq_sstl_in;
	input [1:0]	dqs_diff_in_0;
	input [1:0]	dqs_diff_in_1;
	input [1:0]	dqs_diff_in_2;
	input [1:0]	dqs_diff_in_3;
	input [1:0]	dqs_sstl_n_0;
	input [1:0]	dqs_sstl_n_1;
	input [1:0]	dqs_sstl_n_2;
	input [1:0]	dqs_sstl_n_3;
	input [1:0]	dqs_sstl_p_0;
	input [1:0]	dqs_sstl_p_1;
	input [1:0]	dqs_sstl_p_2;
	input [1:0]	dqs_sstl_p_3;
	input [5:0]	dzoutx;
	input	early_bhniotri;
	input	early_csren;
	input	early_enrnsl;
	input	early_frzreg;
	input	early_nfrzdrv;
	input	early_niotri;
	input	early_plniotri;
	input	early_usrmode;
	input	enrnsl;
	input	entest;
	output [2:0]	fb_clkout;
	input [12*1-1:0]	fr_in_clk;
	input [12*1-1:0]	fr_out_clk;
	input	frzreg;
	output	hps_to_core_ctrl_en;
	input [12*1-1:0]	hr_in_clk;
	input [12*1-1:0]	hr_out_clk;
	input	i50u_ref;
	input	ibp50u;
	input	ibp50u_cal;
	output [5:0]	ioereg_locked;
	input	jtag_clk;
	input	jtag_highz;
	input	jtag_mode;
	input	jtag_sdin;
	output	jtag_sdout;
	input	jtag_shftdr;
	input	jtag_updtdr;
	output	lane_cal_done;
	output	local_bhniotri;
	output	local_enrnsl;
	output	local_frzreg;
	output	local_nfrzdrv;
	output	local_niotri;
	output	local_plniotri;
	output	local_usrmode;
	output	local_wkpullup;
	output [1:0]	lvds_rx_clk_chnl0;
	output [1:0]	lvds_rx_clk_chnl1;
	output [1:0]	lvds_rx_clk_chnl2;
	output [1:0]	lvds_rx_clk_chnl3;
	output [1:0]	lvds_rx_clk_chnl4;
	output [1:0]	lvds_rx_clk_chnl5;
	output [1:0]	lvds_tx_clk_chnl0;
	output [1:0]	lvds_tx_clk_chnl1;
	output [1:0]	lvds_tx_clk_chnl2;
	output [1:0]	lvds_tx_clk_chnl3;
	output [1:0]	lvds_tx_clk_chnl4;
	output [1:0]	lvds_tx_clk_chnl5;
	input [15:0]	mrnk_read_core;
	input [15:0]	mrnk_write_core;
	output [5:0]	n_crnt_clk;
	output [5:0]	n_next_clk;
	input [12*1-1:0]	naclr;
	input [12*1-1:0]	ncein;
	input [12*1-1:0]	nceout;
	output [5:0]	next_clk;
	input	nfrzdrv;
	input	niotri;
	input [12*1-1:0]	nsclr;
	output [11:0]	oct_enable;
	input [47:0]	oeb_from_core;
	input	osc_en_n;
	input	osc_enable_in;
	input	osc_mode_in;
	output	osc_rocount_to_core;
	input	osc_sel_n;
	input [4:0]	phy_clk;
	input [7:0]	phy_clk_phs;
	input	pipeline_global_en_n;
	input	pll_clk;
	input	pll_locked;
	input	plniotri;
	input [12*1-1:0]	progctl;
	input [12*1-1:0]	progoe;
	input [12*1-1:0]	progout;
	input [3:0]	rdata_en_full_core;
	output [3:0]	rdata_valid_core;
	input	regulator_clk;
	input	reinit;
	input	reset_n;
	input	scan_shift_n;
	input [5:0]	scanin;
	output [5:0]	scanout;
	input [5:0]	switch_dn;
	input [5:0]	switch_up;
	input	sync_clk_bot_in;
	output	sync_clk_bot_out;
	input	sync_clk_top_in;
	output	sync_clk_top_out;
	input	sync_data_bot_in;
	output	sync_data_bot_out;
	input	sync_data_top_in;
	output	sync_data_top_out;
	input	test_avl_clk_in_en_n;
	input	test_clk;
	input	test_clk_ph_buf_en_n;
	input	test_clk_pll_en_n;
	input	test_clr_n;
	input	test_datovr_en_n;
	input	test_db_csr_in;
	output [11:0]	test_dbg_in;
	input [11:0]	test_dbg_out;
	input	test_dqs_csr_in;
	input	test_dqs_enable_en_n;
	input	test_fr_clk_en_n;
	input	test_hr_clk_en_n;
	input	test_int_clk_en_n;
	input	test_interp_clk_en_n;
	output	test_ioereg2_csr_out;
	input	test_phy_clk_en_n;
	input	test_phy_clk_lane_en_n;
	input	test_pst_clk_en_n;
	input	test_pst_dll_i;
	output	test_pst_dll_o;
	input	test_tdf_select_n;
	output	test_vref_csr_out;
	output	test_xor_clk;
	input [12*1-1:0]	tpctl;
	output [12*1-1:0]	tpdata;
	input [12*1-1:0]	tpin;
	input [5:0]	up_ph;
	input	usrmode;
	input	vref_ext;
	output	vref_int;
	output [11:0]	weak_pullup_enable;
	input	wkpullup;
	output	x1024_osc_out;
	output	xor_vref;
	input	xprio_clk;
	input	xprio_sync;
	input [7:0]	xprio_xbus;

parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_ac_dqs_dm_dq = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_data_buffer_ctrl = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_db_oe_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_db_out_bypass = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_db_pin_type = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_memory_standard = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_oe_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_rb_sel_ac_hmc_ena = "";
parameter data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_wr_datapath_prgmnvrt = "";
parameter data_buffer__data_buffer_out_if_inst__HIERARCHY = "";
parameter data_buffer__rdwr_buffer_inst_0__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_0__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_0__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_0__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_0__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_0__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_0__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_0__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_1__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_1__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_1__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_1__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_1__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_1__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_1__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_1__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_10__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_10__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_10__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_10__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_10__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_10__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_10__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_10__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_11__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_11__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_11__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_11__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_11__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_11__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_11__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_11__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_2__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_2__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_2__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_2__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_2__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_2__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_2__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_2__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_3__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_3__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_3__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_3__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_3__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_3__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_3__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_3__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_4__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_4__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_4__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_4__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_4__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_4__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_4__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_4__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_5__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_5__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_5__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_5__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_5__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_5__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_5__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_5__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_6__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_6__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_6__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_6__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_6__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_6__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_6__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_6__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_7__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_7__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_7__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_7__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_7__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_7__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_7__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_7__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_8__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_8__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_8__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_8__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_8__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_8__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_8__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_8__a_wr_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_9__a_data_buffer_ctrl = "";
parameter data_buffer__rdwr_buffer_inst_9__a_db_in_bypass = "";
parameter data_buffer__rdwr_buffer_inst_9__a_dbc_sel = "";
parameter data_buffer__rdwr_buffer_inst_9__a_oe_datapath_mod = "";
parameter data_buffer__rdwr_buffer_inst_9__a_pipeline = "";
parameter data_buffer__rdwr_buffer_inst_9__a_prbs = "";
parameter data_buffer__rdwr_buffer_inst_9__a_wdb_bypass = "";
parameter data_buffer__rdwr_buffer_inst_9__a_wr_datapath_mod = "";
parameter data_buffer__HIERARCHY = "";
parameter data_buffer__a_calibration = "";
parameter data_buffer__a_data_buffer_ctrl = "";
parameter data_buffer__a_dft_mode = "";
parameter data_buffer__a_memory_standard = "";
parameter data_buffer__a_mode_rate_in = "";
parameter data_buffer__a_mode_rate_out = "";
parameter [8-1:0] data_buffer__a_phy_wlat = 8'h00;
parameter [8-1:0] data_buffer__a_pipe_latency = 8'h00;
parameter [6-1:0] data_buffer__a_rb_afi_rlat_vlu = 6'b0;
parameter [6-1:0] data_buffer__a_rb_afi_wlat_vlu = 6'b0;
parameter data_buffer__a_rb_avl_ena = "";
parameter data_buffer__a_rb_bc_id_ena = "";
parameter data_buffer__a_rb_burst_length_mode = "";
parameter data_buffer__a_rb_crc_dq0 = "";
parameter data_buffer__a_rb_crc_dq1 = "";
parameter data_buffer__a_rb_crc_dq2 = "";
parameter data_buffer__a_rb_crc_dq3 = "";
parameter data_buffer__a_rb_crc_dq4 = "";
parameter data_buffer__a_rb_crc_dq5 = "";
parameter data_buffer__a_rb_crc_dq6 = "";
parameter data_buffer__a_rb_crc_dq7 = "";
parameter data_buffer__a_rb_crc_dq8 = "";
parameter data_buffer__a_rb_crc_en = "";
parameter data_buffer__a_rb_data_alignment_mode = "";
parameter data_buffer__a_rb_db2core_registered = "";
parameter [4-1:0] data_buffer__a_rb_db_feature = 4'h0;
parameter [7-1:0] data_buffer__a_rb_dbc_wb_reserved_entry = 7'h04;
parameter data_buffer__a_rb_dbi_rd_en = "";
parameter data_buffer__a_rb_dbi_sel = "";
parameter data_buffer__a_rb_dbi_wr_en = "";
parameter data_buffer__a_rb_dft_hmc_phy = "";
parameter data_buffer__a_rb_dft_lbk_phy = "";
parameter data_buffer__a_rb_dft_mux_speed_in = "";
parameter data_buffer__a_rb_dft_mux_speed_out = "";
parameter data_buffer__a_rb_dft_prbs_mode = "";
parameter data_buffer__a_rb_dft_speed_test = "";
parameter data_buffer__a_rb_gpio_0 = "";
parameter data_buffer__a_rb_gpio_1 = "";
parameter data_buffer__a_rb_gpio_10 = "";
parameter data_buffer__a_rb_gpio_11 = "";
parameter data_buffer__a_rb_gpio_2 = "";
parameter data_buffer__a_rb_gpio_3 = "";
parameter data_buffer__a_rb_gpio_4 = "";
parameter data_buffer__a_rb_gpio_5 = "";
parameter data_buffer__a_rb_gpio_6 = "";
parameter data_buffer__a_rb_gpio_7 = "";
parameter data_buffer__a_rb_gpio_8 = "";
parameter data_buffer__a_rb_gpio_9 = "";
parameter data_buffer__a_rb_hmc_or_core = "";
parameter data_buffer__a_rb_mrnk_read_registered = "";
parameter data_buffer__a_rb_mrnk_write_registered = "";
parameter data_buffer__a_rb_phy_clk0_ena = "";
parameter data_buffer__a_rb_phy_clk1_ena = "";
parameter data_buffer__a_rb_preamble_mode = "";
parameter data_buffer__a_rb_ptr_pipeline = "";
parameter data_buffer__a_rb_qr_or_hr = "";
parameter data_buffer__a_rb_rdata_en_full_registered = "";
parameter data_buffer__a_rb_reset_auto_release = "";
parameter data_buffer__a_rb_rwlat_mode = "";
parameter data_buffer__a_rb_sel_core_clk = "";
parameter [3-1:0] data_buffer__a_rb_seq_rd_en_full_pipeline = 3'h0;
parameter [9-1:0] data_buffer__a_rb_tile_id = 9'h00;
parameter data_buffer__a_rb_x4_or_x8_or_x9 = "";
parameter [8-1:0] data_buffer__a_wl_latency = 8'h00;
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_0__gpio_reg__mode = "";
parameter ioereg_top_0___gpio_wrapper_0__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__HIERARCHY = "";
parameter ioereg_top_0___gpio_wrapper_1__gpio_reg__mode = "";
parameter ioereg_top_0___gpio_wrapper_1__HIERARCHY = "";
parameter [12-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_ck_cmd = 12'h000;
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select = "";
parameter [12-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dqss = 12'h000;
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_mode_output = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_in = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_out = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_octrt = "";
parameter [12-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase = 12'h000;
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_pin_usage = "";
parameter [12-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_wl_latency = 10'h000;
parameter [12-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_ck_cmd = 12'h000;
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select = "";
parameter [12-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dqss = 12'h000;
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_mode_output = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_in = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_out = "";
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_octrt = "";
parameter [12-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase = 12'h000;
parameter ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_pin_usage = "";
parameter [12-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_wl_latency = 10'h000;
parameter ioereg_top_0___ioereg_pnr_x2__HIERARCHY = "";
parameter ioereg_top_0___ioereg_pnr_x2__a_ddr2_oeb = "";
parameter ioereg_top_0___ioereg_pnr_x2__a_dpa_enable = "";
parameter [3-1:0] ioereg_top_0___ioereg_pnr_x2__a_lock_speed = 3'h7;
parameter ioereg_top_0___ioereg_pnr_x2__a_power_down = "";
parameter ioereg_top_0___ioereg_pnr_x2__a_power_down_0 = "";
parameter ioereg_top_0___ioereg_pnr_x2__a_power_down_1 = "";
parameter ioereg_top_0___ioereg_pnr_x2__a_power_down_2 = "";
parameter ioereg_top_0___ioereg_pnr_x2__a_sync_control = "";
parameter ioereg_top_0___HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_0__gpio_reg__mode = "";
parameter ioereg_top_1___gpio_wrapper_0__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__HIERARCHY = "";
parameter ioereg_top_1___gpio_wrapper_1__gpio_reg__mode = "";
parameter ioereg_top_1___gpio_wrapper_1__HIERARCHY = "";
parameter [12-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_ck_cmd = 12'h000;
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select = "";
parameter [12-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dqss = 12'h000;
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_mode_output = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_in = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_out = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_octrt = "";
parameter [12-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase = 12'h000;
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_pin_usage = "";
parameter [12-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_wl_latency = 10'h000;
parameter [12-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_ck_cmd = 12'h000;
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select = "";
parameter [12-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dqss = 12'h000;
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_mode_output = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_in = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_out = "";
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_octrt = "";
parameter [12-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase = 12'h000;
parameter ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_pin_usage = "";
parameter [12-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_wl_latency = 10'h000;
parameter ioereg_top_1___ioereg_pnr_x2__HIERARCHY = "";
parameter ioereg_top_1___ioereg_pnr_x2__a_ddr2_oeb = "";
parameter ioereg_top_1___ioereg_pnr_x2__a_dpa_enable = "";
parameter [3-1:0] ioereg_top_1___ioereg_pnr_x2__a_lock_speed = 3'h7;
parameter ioereg_top_1___ioereg_pnr_x2__a_power_down = "";
parameter ioereg_top_1___ioereg_pnr_x2__a_power_down_0 = "";
parameter ioereg_top_1___ioereg_pnr_x2__a_power_down_1 = "";
parameter ioereg_top_1___ioereg_pnr_x2__a_power_down_2 = "";
parameter ioereg_top_1___ioereg_pnr_x2__a_sync_control = "";
parameter ioereg_top_1___HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_0__gpio_reg__mode = "";
parameter ioereg_top_2___gpio_wrapper_0__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__HIERARCHY = "";
parameter ioereg_top_2___gpio_wrapper_1__gpio_reg__mode = "";
parameter ioereg_top_2___gpio_wrapper_1__HIERARCHY = "";
parameter [12-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_ck_cmd = 12'h000;
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select = "";
parameter [12-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dqss = 12'h000;
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_mode_output = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_in = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_out = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_octrt = "";
parameter [12-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase = 12'h000;
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_pin_usage = "";
parameter [12-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_wl_latency = 10'h000;
parameter [12-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_ck_cmd = 12'h000;
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select = "";
parameter [12-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dqss = 12'h000;
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_mode_output = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_in = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_out = "";
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_octrt = "";
parameter [12-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase = 12'h000;
parameter ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_pin_usage = "";
parameter [12-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_wl_latency = 10'h000;
parameter ioereg_top_2___ioereg_pnr_x2__HIERARCHY = "";
parameter ioereg_top_2___ioereg_pnr_x2__a_ddr2_oeb = "";
parameter ioereg_top_2___ioereg_pnr_x2__a_dpa_enable = "";
parameter [3-1:0] ioereg_top_2___ioereg_pnr_x2__a_lock_speed = 3'h7;
parameter ioereg_top_2___ioereg_pnr_x2__a_power_down = "";
parameter ioereg_top_2___ioereg_pnr_x2__a_power_down_0 = "";
parameter ioereg_top_2___ioereg_pnr_x2__a_power_down_1 = "";
parameter ioereg_top_2___ioereg_pnr_x2__a_power_down_2 = "";
parameter ioereg_top_2___ioereg_pnr_x2__a_sync_control = "";
parameter ioereg_top_2___HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_0__gpio_reg__mode = "";
parameter ioereg_top_3___gpio_wrapper_0__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__HIERARCHY = "";
parameter ioereg_top_3___gpio_wrapper_1__gpio_reg__mode = "";
parameter ioereg_top_3___gpio_wrapper_1__HIERARCHY = "";
parameter [12-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_ck_cmd = 12'h000;
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select = "";
parameter [12-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dqss = 12'h000;
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_mode_output = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_in = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_out = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_octrt = "";
parameter [12-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase = 12'h000;
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_pin_usage = "";
parameter [12-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_wl_latency = 10'h000;
parameter [12-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_ck_cmd = 12'h000;
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select = "";
parameter [12-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dqss = 12'h000;
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_mode_output = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_in = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_out = "";
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_octrt = "";
parameter [12-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase = 12'h000;
parameter ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_pin_usage = "";
parameter [12-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_wl_latency = 10'h000;
parameter ioereg_top_3___ioereg_pnr_x2__HIERARCHY = "";
parameter ioereg_top_3___ioereg_pnr_x2__a_ddr2_oeb = "";
parameter ioereg_top_3___ioereg_pnr_x2__a_dpa_enable = "";
parameter [3-1:0] ioereg_top_3___ioereg_pnr_x2__a_lock_speed = 3'h7;
parameter ioereg_top_3___ioereg_pnr_x2__a_power_down = "";
parameter ioereg_top_3___ioereg_pnr_x2__a_power_down_0 = "";
parameter ioereg_top_3___ioereg_pnr_x2__a_power_down_1 = "";
parameter ioereg_top_3___ioereg_pnr_x2__a_power_down_2 = "";
parameter ioereg_top_3___ioereg_pnr_x2__a_sync_control = "";
parameter ioereg_top_3___HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_0__gpio_reg__mode = "";
parameter ioereg_top_4___gpio_wrapper_0__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__HIERARCHY = "";
parameter ioereg_top_4___gpio_wrapper_1__gpio_reg__mode = "";
parameter ioereg_top_4___gpio_wrapper_1__HIERARCHY = "";
parameter [12-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_ck_cmd = 12'h000;
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select = "";
parameter [12-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dqss = 12'h000;
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_mode_output = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_in = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_out = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_octrt = "";
parameter [12-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase = 12'h000;
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_pin_usage = "";
parameter [12-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_wl_latency = 10'h000;
parameter [12-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_ck_cmd = 12'h000;
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select = "";
parameter [12-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dqss = 12'h000;
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_mode_output = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_in = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_out = "";
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_octrt = "";
parameter [12-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase = 12'h000;
parameter ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_pin_usage = "";
parameter [12-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_wl_latency = 10'h000;
parameter ioereg_top_4___ioereg_pnr_x2__HIERARCHY = "";
parameter ioereg_top_4___ioereg_pnr_x2__a_ddr2_oeb = "";
parameter ioereg_top_4___ioereg_pnr_x2__a_dpa_enable = "";
parameter [3-1:0] ioereg_top_4___ioereg_pnr_x2__a_lock_speed = 3'h7;
parameter ioereg_top_4___ioereg_pnr_x2__a_power_down = "";
parameter ioereg_top_4___ioereg_pnr_x2__a_power_down_0 = "";
parameter ioereg_top_4___ioereg_pnr_x2__a_power_down_1 = "";
parameter ioereg_top_4___ioereg_pnr_x2__a_power_down_2 = "";
parameter ioereg_top_4___ioereg_pnr_x2__a_sync_control = "";
parameter ioereg_top_4___HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_0__gpio_reg__mode = "";
parameter ioereg_top_5___gpio_wrapper_0__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__mode = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__mode = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__mode = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__HIERARCHY = "";
parameter ioereg_top_5___gpio_wrapper_1__gpio_reg__mode = "";
parameter ioereg_top_5___gpio_wrapper_1__HIERARCHY = "";
parameter [12-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_ck_cmd = 12'h000;
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select = "";
parameter [12-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dqss = 12'h000;
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_mode_output = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_in = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_mode_rate_out = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_octrt = "";
parameter [12-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase = 12'h000;
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_pin_usage = "";
parameter [12-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_wl_latency = 10'h000;
parameter [12-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_ck_cmd = 12'h000;
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select = "";
parameter [12-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dqss = 12'h000;
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_mode_output = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_in = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_mode_rate_out = "";
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_octrt = "";
parameter [12-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase = 12'h000;
parameter ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_pin_usage = "";
parameter [12-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_struct_gate_delay = 12'h000;
parameter [13-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_time_core_to_codin = 12'h000;
parameter [10-1:0] ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_wl_latency = 10'h000;
parameter ioereg_top_5___ioereg_pnr_x2__HIERARCHY = "";
parameter ioereg_top_5___ioereg_pnr_x2__a_ddr2_oeb = "";
parameter ioereg_top_5___ioereg_pnr_x2__a_dpa_enable = "";
parameter [3-1:0] ioereg_top_5___ioereg_pnr_x2__a_lock_speed = 3'h7;
parameter ioereg_top_5___ioereg_pnr_x2__a_power_down = "";
parameter ioereg_top_5___ioereg_pnr_x2__a_power_down_0 = "";
parameter ioereg_top_5___ioereg_pnr_x2__a_power_down_1 = "";
parameter ioereg_top_5___ioereg_pnr_x2__a_power_down_2 = "";
parameter ioereg_top_5___ioereg_pnr_x2__a_sync_control = "";
parameter ioereg_top_5___HIERARCHY = "";
parameter vref__a_vref_cal = "";
parameter vref__a_vref_enable = "";
parameter vref__a_vref_offset = "";
parameter vref__a_vref_offsetmode = "";
parameter vref__a_vref_range = "";
parameter vref__a_vref_sel = "";
parameter vref__a_vref_val = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_core_dn_prgmnvrt = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_core_up_prgmnvrt = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_core_updnen = "";
parameter [10-1:0] xio_dll_top__xio_dll_pnr__a_rb_ctl_static = 10'h000;
parameter xio_dll_top__xio_dll_pnr__a_rb_ctlsel = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel0 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel1 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel2 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel3 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel4 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel5 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel6 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel7 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel8 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel9 = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dll_en = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_dll_rst_en = "";
parameter [10-1:0] xio_dll_top__xio_dll_pnr__a_rb_dly_pst = 10'h000;
parameter xio_dll_top__xio_dll_pnr__a_rb_dly_pst_en = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_hps_ctrl_en = "";
parameter xio_dll_top__xio_dll_pnr__a_rb_ndllrst_prgmnvrt = "";
parameter [3-1:0] xio_dll_top__xio_dll_pnr__a_rb_new_dll = 3'b000;
parameter xio_dll_top__xio_dll_pnr__powerdown_mode = "";
parameter xio_dll_top__HIERARCHY = "";
parameter xio_dll_top__dll_func_mode = "";
parameter xio_dll_top__powerdown_mode = "";
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_board_delay = 16'h0000;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_broadcast_enable = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_burst_length = "";
parameter [8-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_cas_latency = 8'h00;
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_cmd_latency = 16'h0000;
parameter [7-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_count_threshold = 7'h00;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_ddr4_search = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_en = "";
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_en_latency = 16'h0000;
parameter [6-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_enable_delay = 6'h00;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_select_a = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_select_b = "";
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_shrink_delay = 16'h0000;
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_shrink_gate_delay = 16'h0000;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_enable_b_rank = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_enable_toggler = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_filter_code = "";
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_io_in_delay = 16'h0000;
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_io_out_delay = 16'h0000;
parameter [2-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_kicker_size = 2'h0;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_lock_edge = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_memory_burst_length = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_memory_dqs_type = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_memory_rank_size = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_memory_standard = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_memory_width = "";
parameter [7-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_min_rd_valid_delay = 7'h00;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_mode_rate_in = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_mode_rate_out = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_mrnk_delay = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_multi_rank_enable = "";
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay = 9'h000;
parameter [9-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay = 9'h000;
parameter [10-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay = 10'h000;
parameter [3-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_oct_size = 3'h1;
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_output_phase = 16'h0000;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_pack_mode = "";
parameter [13-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a = 13'h000;
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_adjust = 16'h0000;
parameter [13-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b = 13'h000;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_phy_clk_mode = "";
parameter [8-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_pipe_latency = 8'h00;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_power_down = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_power_down_0 = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_power_down_1 = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_power_down_2 = "";
parameter [4-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_probe_sel = 4'h0;
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_pst_en_shrink = "";
parameter xio_dqs_lgc_top__dqs_lgc_pnr__a_pst_preamble_mode = "";
parameter [10-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a = 10'h000;
parameter [10-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b = 10'h000;
parameter [7-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay = 7'h00;
parameter [8-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay_adjust = 8'h00;
parameter [8-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_rlat = 8'h00;
parameter [7-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_rlat_rd_valid_delay = 7'h00;
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_time_en_full_to_shrunk_a = 16'h0000;
parameter [16-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_time_en_full_to_shrunk_b = 16'h0000;
parameter [4-1:0] xio_dqs_lgc_top__dqs_lgc_pnr__a_track_speed = 4'h0;
parameter xio_dqs_lgc_top__HIERARCHY = "";
parameter [16-1:0] xio_dqs_lgc_top__a_clock_period = 16'h000;
parameter xio_regulator__a_cr_atbsel0 = "";
parameter xio_regulator__a_cr_atbsel1 = "";
parameter xio_regulator__a_cr_atbsel2 = "";
parameter xio_regulator__a_cr_pd = "";
parameter xio_regulator__a_powerdown_mode = "";
parameter HIERARCHY = "";
parameter [16-1:0] a_board_delay = 16'h0000;
parameter a_calibration = "";
parameter [8-1:0] a_cas_latency = 8'h00;
parameter [12-1:0] a_ck_cmd = 12'h000;
parameter [16-1:0] a_clock_period = 16'h000;
parameter [13-1:0] a_cmd_core_to_codin = 13'h000;
parameter [13-1:0] a_cmd_pipe_latency = 13'h000;
parameter [13-1:0] a_dq_read_latency = 13'h000;
parameter [12-1:0] a_dqss = 12'h040;
parameter a_filter_code = "";
parameter [16-1:0] a_io_in_delay = 16'h0000;
parameter [16-1:0] a_io_out_delay = 16'h0000;
parameter a_lane_usage = "";
parameter a_memory_burst_length = "";
parameter a_memory_controller = "";
parameter a_memory_rank_size = "";
parameter a_memory_standard = "";
parameter a_memory_width = "";
parameter a_mode_rate_in = "";
parameter a_mode_rate_out = "";
parameter [16-1:0] a_output_phase = 16'h0000;
parameter a_phy_clk_mode = "";
parameter [8-1:0] a_pipe_latency = 8'h00;
parameter [13-1:0] a_struct_gate_delay = 13'h000;
parameter [8-1:0] a_wl_latency = 8'h00;
parameter powerdown_mode = "";

`ifndef USE_CSR
initial
begin

	i0.xio_dqs_lgc_top.dqs_lgc_pnr.avl_toggler = 1'b0;

	force csr_en = 1'b0;
	force csr_shift_n = 1'b0;

case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[213].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[213].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[213].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[132].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[132].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[132].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[108].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[108].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[108].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[252].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[252].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[252].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_0__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[214].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[214].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[214].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[133].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[133].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[133].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[109].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[109].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[109].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[253].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[253].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[253].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_1__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[223].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[223].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[223].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[142].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[142].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[142].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[118].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[118].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[118].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[262].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[262].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[262].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_10__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[224].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[224].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[224].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[143].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[143].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[143].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[119].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[119].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[119].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[263].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[263].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[263].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_11__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[215].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[215].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[215].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[134].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[134].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[134].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[110].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[110].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[110].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[254].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[254].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[254].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_2__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[216].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[216].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[216].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[135].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[135].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[135].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[111].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[111].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[111].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[255].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[255].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[255].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_3__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[217].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[217].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[217].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[136].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[136].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[136].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[112].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[112].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[112].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[256].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[256].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[256].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_4__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[218].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[218].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[218].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[137].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[137].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[137].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[113].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[113].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[113].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[257].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[257].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[257].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_5__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[219].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[219].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[219].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[138].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[138].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[138].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[114].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[114].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[114].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[258].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[258].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[258].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_6__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[220].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[220].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[220].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[139].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[139].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[139].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[115].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[115].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[115].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[259].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[259].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[259].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_7__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[221].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[221].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[221].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[140].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[140].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[140].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[116].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[116].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[116].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[260].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[260].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[260].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_8__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_ac_dqs_dm_dq)
	"dq_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	"dm_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
	end
	"ac_type" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_db_oe_bypass)
	"db_oe_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[222].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_oe_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[222].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[222].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_db_out_bypass)
	"db_out_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[141].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_out_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[141].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[141].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_oe_datapath_prgmnvrt)
	"oe_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[117].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[117].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[117].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_rb_sel_ac_hmc_ena)
	"sel_ac_hmc_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[261].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel_ac_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[261].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[261].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__data_buffer_out_if_inst__io_data_buffer_out_mux_inst_9__a_wr_datapath_prgmnvrt)
	"wr_datapath_non_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_invert" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_0__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[120].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[120].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[120].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_0__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_0__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_0__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[201].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[201].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[201].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_0__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_0__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_1__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[121].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[121].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[121].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_1__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_1__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_1__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[202].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[202].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[202].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_1__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_1__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_10__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[130].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[130].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[130].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_10__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_10__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[104].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[105].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[104].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[105].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[104].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[105].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_10__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[211].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[211].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[211].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_10__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_10__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_11__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[131].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[131].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[131].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_11__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_11__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[106].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[107].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[106].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[107].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[106].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[107].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_11__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[212].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[212].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[212].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_11__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_11__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_2__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[122].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[122].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[122].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_2__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_2__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_2__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[203].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[203].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[203].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_2__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_2__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_3__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[123].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[123].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[123].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_3__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_3__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_3__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[204].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[204].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[204].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_3__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_3__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_4__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[124].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[124].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[124].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_4__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_4__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_4__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[205].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[205].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[205].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_4__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_4__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_5__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[125].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[125].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[125].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_5__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_5__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_5__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[206].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[206].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[206].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_5__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_5__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_6__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[126].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[126].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[126].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_6__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_6__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_6__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[207].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[207].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[207].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_6__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_6__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_7__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[127].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[127].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[127].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_7__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_7__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_7__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[208].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[208].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[208].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_7__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_7__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_8__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[128].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[128].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[128].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_8__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_8__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_8__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[209].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[209].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[209].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_8__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_8__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_9__a_db_in_bypass)
	"db_in_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[129].csr_reg_bit.csr_reg = 1'b0;
	end
	"db_in_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[129].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[129].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_9__a_dbc_sel)
	"sel_core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_dbc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_9__a_oe_datapath_mod)
	"oe_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[102].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[103].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[102].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[103].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[102].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[103].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_9__a_prbs)
	"sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[210].csr_reg_bit.csr_reg = 1'b1;
	end
	"not_sel_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[210].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[210].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_9__a_wdb_bypass)
	"wdb_not_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
	end
	"wdb_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__rdwr_buffer_inst_9__a_wr_datapath_mod)
	"wr_datapath_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"wr_datapath_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[237].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_rlat_vlu[0];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[238].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_rlat_vlu[1];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[239].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_rlat_vlu[2];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[240].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_rlat_vlu[3];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[241].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_rlat_vlu[4];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[242].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_rlat_vlu[5];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[231].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_wlat_vlu[0];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[232].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_wlat_vlu[1];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[233].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_wlat_vlu[2];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[234].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_wlat_vlu[3];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[235].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_wlat_vlu[4];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[236].csr_reg_bit.csr_reg = data_buffer__a_rb_afi_wlat_vlu[5];
case (data_buffer__a_rb_avl_ena)
	"avl_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[200].csr_reg_bit.csr_reg = 1'b0;
	end
	"avl_enable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[200].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[200].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_bc_id_ena)
	"bc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[162].csr_reg_bit.csr_reg = 1'b0;
	end
	"bc_enable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[162].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[162].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_burst_length_mode)
	"bl8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[276].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[277].csr_reg_bit.csr_reg = 1'b0;
	end
	"bl4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[276].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[277].csr_reg_bit.csr_reg = 1'b0;
	end
	"bl2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[276].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[277].csr_reg_bit.csr_reg = 1'b1;
	end
	"bl_reserved" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[276].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[277].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[276].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[277].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq0)
	"crc_dq0_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq0_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq0_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq0_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq0_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq0_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq0_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq0_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq0_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq0_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq0_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq0_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq1)
	"crc_dq1_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq1_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq1_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq1_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq1_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq1_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq1_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq1_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq1_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq1_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq1_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq1_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq2)
	"crc_dq2_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq2_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq2_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq2_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq2_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq2_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq2_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq2_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq2_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq2_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq2_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq2_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq3)
	"crc_dq3_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq3_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq3_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq3_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq3_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq3_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq3_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq3_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq3_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq3_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq3_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq3_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq4)
	"crc_dq4_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq4_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq4_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq4_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq4_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq4_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq4_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq4_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq4_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq4_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq4_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq4_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq5)
	"crc_dq5_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq5_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq5_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq5_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq5_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq5_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq5_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq5_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq5_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq5_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq5_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq5_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq6)
	"crc_dq6_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq6_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq6_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq6_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq6_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq6_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq6_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq6_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq6_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq6_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq6_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq6_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq7)
	"crc_dq7_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq7_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq7_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq7_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq7_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq7_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq7_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq7_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq7_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq7_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq7_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq7_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_dq8)
	"crc_dq8_pin0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq8_pin1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq8_pin2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq8_pin3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq8_pin4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq8_pin5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq8_pin6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq8_pin7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_dq8_pin8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq8_pin9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq8_pin10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b1;
	end
	"crc_dq8_pin11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_crc_en)
	"crc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[152].csr_reg_bit.csr_reg = 1'b0;
	end
	"crc_en" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[152].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[152].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_data_alignment_mode)
	"align_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[248].csr_reg_bit.csr_reg = 1'b0;
	end
	"align_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[248].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[248].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__a_rb_db2core_registered)
	"not_registered" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[251].csr_reg_bit.csr_reg = 1'b0;
	end
	"registered" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[251].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[251].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[296].csr_reg_bit.csr_reg = data_buffer__a_rb_db_feature[0];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[297].csr_reg_bit.csr_reg = data_buffer__a_rb_db_feature[1];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[298].csr_reg_bit.csr_reg = data_buffer__a_rb_db_feature[2];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[299].csr_reg_bit.csr_reg = data_buffer__a_rb_db_feature[3];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[269].csr_reg_bit.csr_reg = data_buffer__a_rb_dbc_wb_reserved_entry[0];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[270].csr_reg_bit.csr_reg = data_buffer__a_rb_dbc_wb_reserved_entry[1];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[271].csr_reg_bit.csr_reg = data_buffer__a_rb_dbc_wb_reserved_entry[2];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[272].csr_reg_bit.csr_reg = data_buffer__a_rb_dbc_wb_reserved_entry[3];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[273].csr_reg_bit.csr_reg = data_buffer__a_rb_dbc_wb_reserved_entry[4];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[274].csr_reg_bit.csr_reg = data_buffer__a_rb_dbc_wb_reserved_entry[5];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[275].csr_reg_bit.csr_reg = data_buffer__a_rb_dbc_wb_reserved_entry[6];
case (data_buffer__a_rb_dbi_rd_en)
	"dbi_rd_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[268].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_rd_enable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[268].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[268].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_dbi_sel)
	"dbi_dq7" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_dq8" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b1;
	end
	"dbi_dq9" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b1;
	end
	"dbi_dq10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b1;
	end
	"dbi_dq11" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b1;
	end
	"dbi_dq0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_dq1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_dq2" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_dq3" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_dq4" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_dq5" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_dq6" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_dbi_wr_en)
	"dbi_wr_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[149].csr_reg_bit.csr_reg = 1'b0;
	end
	"dbi_wr_enable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[149].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[149].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_dft_hmc_phy)
	"lbk_hmc_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[229].csr_reg_bit.csr_reg = 1'b0;
	end
	"lbk_hmc_enable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[229].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[229].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_dft_lbk_phy)
	"lbk_phy_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[228].csr_reg_bit.csr_reg = 1'b0;
	end
	"lbk_phy_enable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[228].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[228].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_dft_mux_speed_in)
	"sel_speed_in0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[265].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_speed_in1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[265].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[265].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_dft_mux_speed_out)
	"sel_speed_out0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[266].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_speed_out1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[266].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[266].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_dft_prbs_mode)
	"oe_0_dq_0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_0_dq_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_1_dq_0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_1_dq_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b0;
	end
	"oe_prbs_dq_0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b1;
	end
	"oe_prbs_dq_prbs" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b1;
	end
	"oe_0_dq_01" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b1;
	end
	"oe_0_dq_10" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_dft_speed_test)
	"sel_speed_test_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[267].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel_speed_test_enable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[267].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[267].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_0)
	"gpio_0_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[281].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_0_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[281].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[281].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_1)
	"gpio_1_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[282].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_1_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[282].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[282].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_10)
	"gpio_10_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[291].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_10_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[291].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[291].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_11)
	"gpio_11_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[292].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_11_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[292].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[292].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_2)
	"gpio_2_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[283].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_2_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[283].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[283].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_3)
	"gpio_3_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[284].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_3_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[284].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[284].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_4)
	"gpio_4_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[285].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_4_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[285].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[285].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_5)
	"gpio_5_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[286].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_5_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[286].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[286].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_6)
	"gpio_6_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[287].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_6_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[287].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[287].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_7)
	"gpio_7_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[288].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_7_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[288].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[288].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_8)
	"gpio_8_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[289].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_8_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[289].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[289].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_gpio_9)
	"gpio_9_false" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[290].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_9_true" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[290].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[290].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_hmc_or_core)
	"core" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[144].csr_reg_bit.csr_reg = 1'b0;
	end
	"hmc" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[144].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[144].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_mrnk_read_registered)
	"mrnk_read_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[279].csr_reg_bit.csr_reg = 1'b0;
	end
	"mrnk_read_registered" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[279].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[279].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_mrnk_write_registered)
	"mrnk_write_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[280].csr_reg_bit.csr_reg = 1'b0;
	end
	"mrnk_write_registered" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[280].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[280].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_phy_clk0_ena)
	"phy_clk0_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[249].csr_reg_bit.csr_reg = 1'b0;
	end
	"phy_clk0_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[249].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[249].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__a_rb_phy_clk1_ena)
	"phy_clk1_disable" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[250].csr_reg_bit.csr_reg = 1'b0;
	end
	"phy_clk1_ena" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[250].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[250].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__a_rb_preamble_mode)
	"preamble_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[246].csr_reg_bit.csr_reg = 1'b0;
	end
	"preamble_two_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[246].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[246].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_ptr_pipeline)
	"ptr_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[243].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[244].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[245].csr_reg_bit.csr_reg = 1'b0;
	end
	"ptr_one_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[243].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[244].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[245].csr_reg_bit.csr_reg = 1'b0;
	end
	"ptr_two_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[243].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[244].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[245].csr_reg_bit.csr_reg = 1'b0;
	end
	"ptr_three_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[243].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[244].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[245].csr_reg_bit.csr_reg = 1'b0;
	end
	"ptr_four_cycle" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[243].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[244].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[245].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[243].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[244].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[245].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_qr_or_hr)
	"hr" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[199].csr_reg_bit.csr_reg = 1'b0;
	end
	"qr" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[199].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[199].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_rdata_en_full_registered)
	"rdata_en_full_bypass" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[278].csr_reg_bit.csr_reg = 1'b0;
	end
	"rdata_en_full_registered" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[278].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[278].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_reset_auto_release)
	"avl_release" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[247].csr_reg_bit.csr_reg = 1'b0;
	end
	"auto_release" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[247].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[247].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (data_buffer__a_rb_rwlat_mode)
	"csr_vlu" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[230].csr_reg_bit.csr_reg = 1'b0;
	end
	"avl_vlu" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[230].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[230].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (data_buffer__a_rb_sel_core_clk)
	"phy_clk0" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[264].csr_reg_bit.csr_reg = 1'b0;
	end
	"phy_clk1" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[264].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[264].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[293].csr_reg_bit.csr_reg = data_buffer__a_rb_seq_rd_en_full_pipeline[0];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[294].csr_reg_bit.csr_reg = data_buffer__a_rb_seq_rd_en_full_pipeline[1];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[295].csr_reg_bit.csr_reg = data_buffer__a_rb_seq_rd_en_full_pipeline[2];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[153].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[0];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[154].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[1];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[155].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[2];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[156].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[3];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[157].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[4];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[158].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[5];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[159].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[6];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[160].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[7];
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[161].csr_reg_bit.csr_reg = data_buffer__a_rb_tile_id[8];
case (data_buffer__a_rb_x4_or_x8_or_x9)
	"x9_mode" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[150].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[151].csr_reg_bit.csr_reg = 1'b0;
	end
	"x8_mode" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[150].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[151].csr_reg_bit.csr_reg = 1'b0;
	end
	"x4_mode" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[150].csr_reg_bit.csr_reg = 1'b0;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[151].csr_reg_bit.csr_reg = 1'b1;
	end
	"reserved" : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[150].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[151].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[150].csr_reg_bit.csr_reg = 1'b1;
		force i0.data_buffer.data_buffer_cnfg_inst.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[151].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[0];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[1];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[10];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[11];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[2];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[3];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[4];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[5];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[6];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[7];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[8];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[9];
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[0];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[1];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[10];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[11];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[2];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[3];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[4];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[5];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[6];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[7];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[8];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[9];
case (ioereg_top_0___ioereg_pnr_x2__a_ddr2_oeb)
	"ddr3_preamble" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"ddr2_preamble" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__a_dpa_enable)
	"dpa_disabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"dpa_enabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__a_lock_speed[0];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__a_lock_speed[1];
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = ioereg_top_0___ioereg_pnr_x2__a_lock_speed[2];
case (ioereg_top_0___ioereg_pnr_x2__a_power_down)
	"power_on" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__a_power_down_0)
	"power_on_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_0" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__a_power_down_1)
	"power_on_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_1" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__a_power_down_2)
	"power_on_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_2" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_0___ioereg_pnr_x2__a_sync_control)
	"sync_disabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"sync_enabled" : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_0_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[0];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[1];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[10];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[11];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[2];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[3];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[4];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[5];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[6];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[7];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[8];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[9];
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[0];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[1];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[10];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[11];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[2];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[3];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[4];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[5];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[6];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[7];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[8];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[9];
case (ioereg_top_1___ioereg_pnr_x2__a_ddr2_oeb)
	"ddr3_preamble" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"ddr2_preamble" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__a_dpa_enable)
	"dpa_disabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"dpa_enabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__a_lock_speed[0];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__a_lock_speed[1];
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = ioereg_top_1___ioereg_pnr_x2__a_lock_speed[2];
case (ioereg_top_1___ioereg_pnr_x2__a_power_down)
	"power_on" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__a_power_down_0)
	"power_on_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_0" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__a_power_down_1)
	"power_on_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_1" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__a_power_down_2)
	"power_on_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_2" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_1___ioereg_pnr_x2__a_sync_control)
	"sync_disabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"sync_enabled" : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_1_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[0];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[1];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[10];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[11];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[2];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[3];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[4];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[5];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[6];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[7];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[8];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[9];
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[0];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[1];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[10];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[11];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[2];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[3];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[4];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[5];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[6];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[7];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[8];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[9];
case (ioereg_top_2___ioereg_pnr_x2__a_ddr2_oeb)
	"ddr3_preamble" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"ddr2_preamble" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__a_dpa_enable)
	"dpa_disabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"dpa_enabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__a_lock_speed[0];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__a_lock_speed[1];
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = ioereg_top_2___ioereg_pnr_x2__a_lock_speed[2];
case (ioereg_top_2___ioereg_pnr_x2__a_power_down)
	"power_on" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__a_power_down_0)
	"power_on_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_0" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__a_power_down_1)
	"power_on_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_1" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__a_power_down_2)
	"power_on_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_2" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_2___ioereg_pnr_x2__a_sync_control)
	"sync_disabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"sync_enabled" : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_2_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[0];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[1];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[10];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[11];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[2];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[3];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[4];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[5];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[6];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[7];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[8];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[9];
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[0];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[1];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[10];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[11];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[2];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[3];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[4];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[5];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[6];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[7];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[8];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[9];
case (ioereg_top_3___ioereg_pnr_x2__a_ddr2_oeb)
	"ddr3_preamble" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"ddr2_preamble" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__a_dpa_enable)
	"dpa_disabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"dpa_enabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__a_lock_speed[0];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__a_lock_speed[1];
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = ioereg_top_3___ioereg_pnr_x2__a_lock_speed[2];
case (ioereg_top_3___ioereg_pnr_x2__a_power_down)
	"power_on" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__a_power_down_0)
	"power_on_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_0" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__a_power_down_1)
	"power_on_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_1" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__a_power_down_2)
	"power_on_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_2" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_3___ioereg_pnr_x2__a_sync_control)
	"sync_disabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"sync_enabled" : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_3_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[0];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[1];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[10];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[11];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[2];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[3];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[4];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[5];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[6];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[7];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[8];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[9];
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[0];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[1];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[10];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[11];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[2];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[3];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[4];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[5];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[6];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[7];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[8];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[9];
case (ioereg_top_4___ioereg_pnr_x2__a_ddr2_oeb)
	"ddr3_preamble" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"ddr2_preamble" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__a_dpa_enable)
	"dpa_disabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"dpa_enabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__a_lock_speed[0];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__a_lock_speed[1];
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = ioereg_top_4___ioereg_pnr_x2__a_lock_speed[2];
case (ioereg_top_4___ioereg_pnr_x2__a_power_down)
	"power_on" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__a_power_down_0)
	"power_on_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_0" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__a_power_down_1)
	"power_on_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_1" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__a_power_down_2)
	"power_on_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_2" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_4___ioereg_pnr_x2__a_sync_control)
	"sync_disabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"sync_enabled" : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_4_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_0__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xin_dlychn0__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xin_dlychn1__a_rb_ireg_dlychn_sel)
	"dly_setting_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_9" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_10" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_11" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_12" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_13" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_14" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_15" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_16" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_17" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_18" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_19" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_20" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_21" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_22" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_23" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_24" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_25" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_26" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_27" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_28" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_29" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_30" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_31" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_32" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_33" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_34" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_35" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_36" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_37" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_38" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_39" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_40" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_41" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_42" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_43" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_44" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_45" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_46" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_47" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_48" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_4" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_49" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_50" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_51" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_52" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_53" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_54" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_55" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_56" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_57" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_58" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_5" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_59" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_60" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_61" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_62" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_63" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b1;
	end
	"dly_setting_6" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_7" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_setting_8" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_fr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_fr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_hr_in_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_hr_out_clk__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_iodout0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_iodout1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_iodout2__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_iodout3__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_naclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_ncein__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_nceout__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_noe0__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_noe1__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xinv_nsclr__a_rb_sel)
	"in_buf" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"in_inv" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_dfm__a_rb_ireg_or_oreg_sel)
	"outreg_input" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
	end
	"buffer_input" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_halfrate_oreg_ereg__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_fr_out_clk_ereg_ena)
	"fr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_hr_out_clk_ereg_ena)
	"hr_out_clk_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_out_clk_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_ena)
	"naclr_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_naclr_ereg_sel)
	"ereg_nclr_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_npre_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nceout_ereg_ena)
	"nceout_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_clk_rst_gen__a_rb_nsclr_ereg_ena)
	"nsclr_ereg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ereg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__xio_gpio_oe_reg__a_rb_ereg_sclr_val)
	"ereg_sclr_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_sclr_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ereg__a_rb_ereg_tieoff_val)
	"ereg_tieoff_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	"ereg_tieoff_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux0__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux1__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux2__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_4to1_mux3__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_ddio_in__a_rb_sclr_val)
	"sclr_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	"sclr_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_fr_in_clk_ena)
	"fr_in_clk_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	"fr_in_clk_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_hr_in_clk_ena)
	"hr_in_clk_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b1;
	end
	"hr_in_clk_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_ena)
	"naclr_ireg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_ireg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_naclr_ireg_sel)
	"ireg_nclr_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	"ireg_npre_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_ncein_ireg_ena)
	"ncein_ireg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	"ncein_ireg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_ireg__xio_gpio_in_clk_rst_gen__a_rb_nsclr_ireg_ena)
	"nsclr_ireg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_ireg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oe_dly_chn__a_rb_ereg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_4to1_mux__a_rb_mux_sel)
	"sel0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	"sel2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	"sel3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_ddr_ena)
	"oreg_ddr_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_ddr_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_ddio_out__a_rb_oreg_sclr_val)
	"oreg_sclr_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_sclr_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_0__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_halfrate_oreg_ereg_1__a_rb_hr_reg_byp)
	"hr_reg_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_reg_bypass_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_fr_out_clk_oreg_ena)
	"fr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
	end
	"fr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_hr_out_clk_oreg_ena)
	"hr_out_clk_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"hr_out_clk_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_ena)
	"naclr_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	"naclr_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_naclr_oreg_sel)
	"oreg_nclr_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_npre_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nceout_oreg_ena)
	"nceout_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"nceout_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__xio_gpio_out_clk_rst_gen__a_rb_nsclr_oreg_ena)
	"nsclr_oreg_dis" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"nsclr_oreg_ena" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_oreg__a_rb_oreg_tieoff_val)
	"oreg_tieoff_val_low" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"oreg_tieoff_val_high" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_gpio_out_dly_chn__a_rb_oreg_dlychn_sel)
	"outdly_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_9" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_10" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_11" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_12" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_13" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_14" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_15" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"outdly_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_3" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_4" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_5" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_6" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_7" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"outdly_8" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_debug)
	"jtag_debug_off" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_debug_on" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_din_or_pll_sel)
	"jtag_din_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_pll_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___gpio_wrapper_1__gpio_reg__xio_jtag__a_rb_gpio_or_ddr_sel)
	"jtag_gpio_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"jtag_ddr_sel" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[0];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[1];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[10];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[11];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[2];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[3];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[4];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[5];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[6];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[7];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[8];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_0.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_0__a_output_phase[9];
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dfx_mode)
	"dfx_disabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_mcu_probe" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	"dfx_dqs_gate_probe" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	"dfx_dq_dqs_probe" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dq_select)
	"dq_disabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_sstl_in" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_loopback_in" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_xor_loopback_in" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	"dq_differential_in" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_out" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_x12_out" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	"dq_differential_in_avl_x12_out" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dqs_select)
	"dqs_sampler_b_a_rise" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_fall" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_a" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_sampler_b_a_over" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_over" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_b_a_rank" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	"dqs_sampler_a_b_rank" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_dynoct)
	"oct_enabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	"oct_disabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_gpio_differential)
	"gpio_single_ended" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	"gpio_differential" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_initial_out)
	"initial_out_z" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	"initial_out_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	"initial_out_x" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b1;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = 1'b0;
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_mode_ddr)
	"mode_sdr" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b0;
	end
	"mode_ddr" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_octrt)
	"static_oct_off" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	"static_oct_on" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[0];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[1];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[10];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[11];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[2];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[3];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[4];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[5];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[6];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[7];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[8];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_pnr_1.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__ioereg_pnr_1__a_output_phase[9];
case (ioereg_top_5___ioereg_pnr_x2__a_ddr2_oeb)
	"ddr3_preamble" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	"ddr2_preamble" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__a_dpa_enable)
	"dpa_disabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"dpa_enabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__a_lock_speed[0];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__a_lock_speed[1];
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = ioereg_top_5___ioereg_pnr_x2__a_lock_speed[2];
case (ioereg_top_5___ioereg_pnr_x2__a_power_down)
	"power_on" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__a_power_down_0)
	"power_on_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_0" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__a_power_down_1)
	"power_on_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_1" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__a_power_down_2)
	"power_on_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_2" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (ioereg_top_5___ioereg_pnr_x2__a_sync_control)
	"sync_disabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"sync_enabled" : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.ioereg_top_5_.ioereg_pnr_x2.ioereg_misc.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (vref__a_vref_cal)
	"a_vref_cal_enable" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_cal_disable" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (vref__a_vref_enable)
	"a_vref_disable" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_enable" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (vref__a_vref_offset)
	"a_vref_offset_0" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_offset_1" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_offset_2" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_offset_3" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_offset_4" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_offset_5" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_offset_6" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_offset_7" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (vref__a_vref_offsetmode)
	"a_vref_offsetmode_add" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_offsetmode_minus" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (vref__a_vref_range)
	"a_vref_range1" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_range2" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (vref__a_vref_sel)
	"a_vref_sel_ext" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_sel_int" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_sel_loop1" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_sel_byp" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_sel_loop2" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (vref__a_vref_val)
	"a_vref_val_0" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_1" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_2" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_3" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_4" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_5" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_6" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_7" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_8" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_9" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_10" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_11" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_12" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_13" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_14" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_15" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_16" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_17" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_18" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_19" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_20" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_21" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_22" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_23" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_24" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_25" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_26" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_27" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_28" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_29" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_30" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_31" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_vref_val_32" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_33" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_34" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_35" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_36" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_37" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_38" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_39" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_40" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_41" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_42" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_43" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_44" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_45" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_46" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_47" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_48" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_49" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_vref_val_50" : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.vref.xcsr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_core_dn_prgmnvrt)
	"off" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	"on" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_core_up_prgmnvrt)
	"on" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	"off" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_core_updnen)
	"core_updn_dis" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	"core_updn_en" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[0];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[1];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[2];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[3];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[4];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[5];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[6];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[7];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[8];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_ctl_static[9];
case (xio_dll_top__xio_dll_pnr__a_rb_ctlsel)
	"ctl_dynamic" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
	end
	"ctl_static" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel0)
	"pvt_gry_0" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_0" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_0" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	"dft_dll_reset" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel1)
	"pvt_gry_1" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_1" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_1" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
	end
	"dft_overflow" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel2)
	"pvt_gry_2" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_2" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_2" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"gate_state_0" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel3)
	"pvt_gry_3" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_3" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_3" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
	end
	"gate_state_1" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel4)
	"pvt_gry_4" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_4" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_4" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	"gate_state_2" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel5)
	"pvt_gry_5" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_5" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_5" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	"gate_state_3" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel6)
	"pvt_gry_6" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_6" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_6" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	"gate_state_4" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel7)
	"pvt_gry_7" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_7" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_7" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	"dft_unused1" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel8)
	"pvt_gry_8" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_8" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_8" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
	end
	"dft_unused2" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dftmuxsel9)
	"pvt_gry_9" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
	end
	"pvt_binary_9" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
	end
	"int_binary_9" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
	end
	"dft_ctrl_to_core" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dll_en)
	"dll_dis" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"dll_en" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_dll_rst_en)
	"dll_rst_dis" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"dll_rst_en" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[0];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[1];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[2];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[3];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[4];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[5];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[6];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[7];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[8];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_dly_pst[9];
case (xio_dll_top__xio_dll_pnr__a_rb_dly_pst_en)
	"dly_adj_dis" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	"dly_adj_en" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_hps_ctrl_en)
	"hps_ctrl_dis" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs_2.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"hps_ctrl_en" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs_2.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs_2.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dll_top__xio_dll_pnr__a_rb_ndllrst_prgmnvrt)
	"off" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"on" : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_new_dll[0];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_new_dll[1];
		force i0.xio_dll_top.xio_dll_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = xio_dll_top__xio_dll_pnr__a_rb_new_dll[2];
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_broadcast_enable)
	"disable_broadcast" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"generate_broadcast" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	"top_in_broadcast" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	"bottom_in_broadcast" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[28].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[29].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_burst_length)
	"burst_length_10" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	"burst_length_8" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b1;
	end
	"burst_length_4" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	"burst_length_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[13].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[14].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_count_threshold[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_count_threshold[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_count_threshold[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[4].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_count_threshold[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[5].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_count_threshold[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[6].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_count_threshold[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[7].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_count_threshold[6];
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_ddr4_search)
	"ddr3_search" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	"ddr4_search" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[8].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_en)
	"dqs_gated" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[223].csr_reg_bit.csr_reg = 1'b0;
	end
	"dqs_pass" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[223].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[223].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[15].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_enable_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[16].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_enable_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[17].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_enable_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[18].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_enable_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[19].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_enable_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[20].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_enable_delay[5];
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_select_a)
	"a_dqs_diff_in_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_dqs_diff_in_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_dqs_diff_in_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_dqs_diff_in_3" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_dqs_sstl_p_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_dqs_sstl_p_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_dqs_sstl_p_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_dqs_sstl_p_3" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	"a_dqs_sstl_n_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_dqs_sstl_n_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_dqs_sstl_n_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_dqs_sstl_n_3" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_dqs_loop_back0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_dqs_loop_back1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_constant" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	"a_dqs_interpolator" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[72].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[73].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[74].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[75].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_dqs_select_b)
	"b_dqs_diff_in_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"b_dqs_diff_in_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"b_dqs_diff_in_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"b_dqs_diff_in_3" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"b_dqs_sstl_p_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"b_dqs_sstl_p_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"b_dqs_sstl_p_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"b_dqs_sstl_p_3" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	"b_dqs_sstl_n_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	"b_dqs_sstl_n_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	"b_dqs_sstl_n_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	"b_dqs_sstl_n_3" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	"b_dqs_loop_back0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	"b_dqs_loop_back1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	"b_constant" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	"b_dqs_interpolator" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[76].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[77].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[78].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[79].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_enable_b_rank)
	"disable_b_rank" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[224].csr_reg_bit.csr_reg = 1'b0;
	end
	"enable_b_rank" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[224].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[224].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_enable_toggler)
	"preamble_track_dqs_enable" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = 1'b0;
	end
	"preamble_track_toggler" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[80].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_filter_code)
	"freq_08ghz" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
	end
	"freq_10ghz" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b1;
	end
	"freq_12ghz" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	"freq_16ghz" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[30].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[31].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[39].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_kicker_size[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[40].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_kicker_size[1];
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_lock_edge)
	"preamble_lock_rising_edge" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	"preamble_lock_falling_edge" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_mode_rate_in)
	"in_rate_full" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"in_rate_1_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b1;
	end
	"in_rate_1_4" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[9].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[10].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_mode_rate_out)
	"out_rate_full" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	"out_rate_1_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	"out_rate_1_4" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	"out_rate_1_8" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[11].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[12].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_mrnk_delay)
	"mrnk_short" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[229].csr_reg_bit.csr_reg = 1'b0;
	end
	"mrnk_long" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[229].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[229].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[201].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[202].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[203].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[204].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[205].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[206].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[207].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[208].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[209].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_0_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[120].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[121].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[122].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[123].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[124].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[125].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[126].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[127].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[128].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_10_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[111].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[112].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[113].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[114].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[115].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[116].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[117].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[118].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[119].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_11_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[210].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[211].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[212].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[213].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[214].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[215].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[216].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[217].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[218].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_1_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[192].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[193].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[194].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[195].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[196].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[197].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[198].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[199].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[200].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_2_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[183].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[184].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[185].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[186].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[187].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[188].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[189].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[190].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[191].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_3_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[174].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[175].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[176].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[177].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[178].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[179].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[180].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[181].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[182].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_4_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[165].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[166].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[167].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[168].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[169].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[170].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[171].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[172].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[173].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_5_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[156].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[157].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[158].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[159].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[160].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[161].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[162].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[163].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[164].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_6_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[147].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[148].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[149].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[150].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[151].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[152].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[153].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[154].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[155].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_7_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[138].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[139].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[140].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[141].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[142].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[143].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[144].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[145].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[146].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_8_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[129].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[130].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[131].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[132].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[133].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[134].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[135].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[136].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[137].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dq_9_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[101].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[102].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[103].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[104].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[105].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[106].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[107].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[108].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[109].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[110].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_non_pvt_dqs_delay[9];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[42].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_oct_size[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[43].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_oct_size[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[44].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_oct_size[2];
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_pack_mode)
	"packed" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	"not_packed" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[41].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[46].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[47].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[56].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[10];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[57].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[11];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[58].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[12];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[48].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[49].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[50].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[51].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[52].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[53].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[54].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[55].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_a[9];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[59].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[60].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[69].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[10];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[70].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[11];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[71].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[12];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[61].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[62].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[63].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[64].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[65].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[66].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[67].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[68].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_phase_shift_b[9];
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_phy_clk_mode)
	"phy_clk_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
	end
	"phy_clk_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[45].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_power_down)
	"power_on" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[228].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[228].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[228].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_power_down_0)
	"power_on_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[225].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_power_down_1)
	"power_on_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[226].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_power_down_2)
	"power_on_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b0;
	end
	"power_off_2" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[227].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[219].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_probe_sel[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[220].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_probe_sel[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[221].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_probe_sel[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[222].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_probe_sel[3];
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_pst_en_shrink)
	"shrink_0_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"shrink_0_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b0;
	end
	"shrink_1_0" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	"shrink_1_1" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b1;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[32].csr_reg_bit.csr_reg = 1'b0;
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[33].csr_reg_bit.csr_reg = 1'b1;
	end
	endcase
case (xio_dqs_lgc_top__dqs_lgc_pnr__a_pst_preamble_mode)
	"ddr3_preamble" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	"ddr4_preamble" : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[34].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[91].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[92].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[93].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[94].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[95].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[96].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[97].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[98].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[99].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[100].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_a[9];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[81].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[82].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[83].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[84].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[85].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[86].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[87].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[88].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[7];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[89].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[8];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[90].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_pvt_input_delay_b[9];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[21].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[22].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[23].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[24].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay[3];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[25].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay[4];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[26].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay[5];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[27].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_rd_valid_delay[6];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[35].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_track_speed[0];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[36].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_track_speed[1];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[37].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_track_speed[2];
		force i0.xio_dqs_lgc_top.dqs_lgc_pnr.csr_reg_nregs.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[38].csr_reg_bit.csr_reg = xio_dqs_lgc_top__dqs_lgc_pnr__a_track_speed[3];
case (xio_regulator__a_cr_atbsel0)
	"cr_atbsel0_dis" : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	"cr_atbsel0_en" : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[1].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_regulator__a_cr_atbsel1)
	"cr_atbsel1_dis" : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	"cr_atbsel1_en" : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[2].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_regulator__a_cr_atbsel2)
	"cr_atbsel2_en" : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b1;
	end
	"cr_atbsel2_dis" : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	default : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[3].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase
case (xio_regulator__a_cr_pd)
	"cr_pd_dis" : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	"cr_pd_en" : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b1;
	end
	default : begin
		force i0.xio_regulator.xio_vreg_cnfg.csr_reg_nregs[0].csr_reg_nbits.csr_reg_bit[0].csr_reg_bit.csr_reg = 1'b0;
	end
	endcase

	#111
	force csr_en = 1'b1;
	force csr_shift_n = 1'b1;
end
`endif

io_12_lane__nf5es_abphy i0 (
	.ac_hmc( ac_hmc),
	.afi_rlat_core( afi_rlat_core),
	.afi_wlat_core( afi_wlat_core),
	.atbi_0( atbi_0),
	.atbi_1( atbi_1),
	.atpg_en_n( atpg_en_n),
	.avl_address_in( avl_address_in),
	.avl_address_out( avl_address_out),
	.avl_clk_in( avl_clk_in),
	.avl_clk_out( avl_clk_out),
	.avl_read_in( avl_read_in),
	.avl_read_out( avl_read_out),
	.avl_readdata_in( avl_readdata_in),
	.avl_readdata_out( avl_readdata_out),
	.avl_write_in( avl_write_in),
	.avl_write_out( avl_write_out),
	.avl_writedata_in( avl_writedata_in),
	.avl_writedata_out( avl_writedata_out),
	.bhniotri( bhniotri),
	.broadcast_in_bot( broadcast_in_bot),
	.broadcast_in_top( broadcast_in_top),
	.broadcast_out_bot( broadcast_out_bot),
	.broadcast_out_top( broadcast_out_top),
	.cas_csrdin( cas_csrdin),
	.cas_csrdout( cas_csrdout),
	.cfg_cmd_rate( cfg_cmd_rate),
	.cfg_dbc_ctrl_sel( cfg_dbc_ctrl_sel),
	.cfg_dbc_dualport_en( cfg_dbc_dualport_en),
	.cfg_dbc_in_protocol( cfg_dbc_in_protocol),
	.cfg_dbc_pipe_lat( cfg_dbc_pipe_lat),
	.cfg_dbc_rc_en( cfg_dbc_rc_en),
	.cfg_dbc_slot_offset( cfg_dbc_slot_offset),
	.cfg_dbc_slot_rotate_en( cfg_dbc_slot_rotate_en),
	.cfg_output_regd( cfg_output_regd),
	.cfg_reorder_rdata( cfg_reorder_rdata),
	.cfg_rmw_en( cfg_rmw_en),
	.clk_pll( clk_pll),
	.codin_n( codin_n),
	.codin_nb( codin_nb),
	.codin_p( codin_p),
	.codin_pb( codin_pb),
	.core2dbc_rd_data_rdy( core2dbc_rd_data_rdy),
	.core2dbc_wr_data_vld0( core2dbc_wr_data_vld0),
	.core2dbc_wr_data_vld1( core2dbc_wr_data_vld1),
	.core2dbc_wr_ecc_info( core2dbc_wr_ecc_info),
	.core_dll( core_dll),
	.crnt_clk( crnt_clk),
	.csr_clk( csr_clk),
	.csr_clk_left( csr_clk_left),
	.csr_en( csr_en),
	.csr_en_left( csr_en_left),
	.csr_in( csr_in),
	.csr_out( csr_out),
	.csr_shift_n( csr_shift_n),
	.ctl2dbc_cs0( ctl2dbc_cs0),
	.ctl2dbc_cs1( ctl2dbc_cs1),
	.ctl2dbc_mask_entry0( ctl2dbc_mask_entry0),
	.ctl2dbc_mask_entry1( ctl2dbc_mask_entry1),
	.ctl2dbc_misc0( ctl2dbc_misc0),
	.ctl2dbc_misc1( ctl2dbc_misc1),
	.ctl2dbc_mrnk_read0( ctl2dbc_mrnk_read0),
	.ctl2dbc_mrnk_read1( ctl2dbc_mrnk_read1),
	.ctl2dbc_nop0( ctl2dbc_nop0),
	.ctl2dbc_nop1( ctl2dbc_nop1),
	.ctl2dbc_rb_rdptr0( ctl2dbc_rb_rdptr0),
	.ctl2dbc_rb_rdptr1( ctl2dbc_rb_rdptr1),
	.ctl2dbc_rb_rdptr_vld0( ctl2dbc_rb_rdptr_vld0),
	.ctl2dbc_rb_rdptr_vld1( ctl2dbc_rb_rdptr_vld1),
	.ctl2dbc_rb_wrptr0( ctl2dbc_rb_wrptr0),
	.ctl2dbc_rb_wrptr1( ctl2dbc_rb_wrptr1),
	.ctl2dbc_rb_wrptr_vld0( ctl2dbc_rb_wrptr_vld0),
	.ctl2dbc_rb_wrptr_vld1( ctl2dbc_rb_wrptr_vld1),
	.ctl2dbc_rd_type0( ctl2dbc_rd_type0),
	.ctl2dbc_rd_type1( ctl2dbc_rd_type1),
	.ctl2dbc_rdata_en_full0( ctl2dbc_rdata_en_full0),
	.ctl2dbc_rdata_en_full1( ctl2dbc_rdata_en_full1),
	.ctl2dbc_seq_en0( ctl2dbc_seq_en0),
	.ctl2dbc_seq_en1( ctl2dbc_seq_en1),
	.ctl2dbc_wb_rdptr0( ctl2dbc_wb_rdptr0),
	.ctl2dbc_wb_rdptr1( ctl2dbc_wb_rdptr1),
	.ctl2dbc_wb_rdptr_vld0( ctl2dbc_wb_rdptr_vld0),
	.ctl2dbc_wb_rdptr_vld1( ctl2dbc_wb_rdptr_vld1),
	.ctl2dbc_wrdata_vld0( ctl2dbc_wrdata_vld0),
	.ctl2dbc_wrdata_vld1( ctl2dbc_wrdata_vld1),
	.data_from_core( data_from_core),
	.data_to_core( data_to_core),
	.dbc2core_rd_data_vld0( dbc2core_rd_data_vld0),
	.dbc2core_rd_data_vld1( dbc2core_rd_data_vld1),
	.dbc2core_rd_type( dbc2core_rd_type),
	.dbc2core_wb_pointer( dbc2core_wb_pointer),
	.dbc2core_wr_data_rdy( dbc2core_wr_data_rdy),
	.dbc2ctl_all_rd_done( dbc2ctl_all_rd_done),
	.dbc2ctl_rb_retire_ptr( dbc2ctl_rb_retire_ptr),
	.dbc2ctl_rb_retire_ptr_vld( dbc2ctl_rb_retire_ptr_vld),
	.dbc2ctl_rd_data_vld( dbc2ctl_rd_data_vld),
	.dbc2ctl_wb_retire_ptr( dbc2ctl_wb_retire_ptr),
	.dbc2ctl_wb_retire_ptr_vld( dbc2ctl_wb_retire_ptr_vld),
	.dbc2db_wb_wrptr( dbc2db_wb_wrptr),
	.dbc2db_wb_wrptr_vld( dbc2db_wb_wrptr_vld),
	.dft_core2db( dft_core2db),
	.dft_db2core( dft_db2core),
	.dft_phy_clk( dft_phy_clk),
	.dft_prbs_done( dft_prbs_done),
	.dft_prbs_ena_n( dft_prbs_ena_n),
	.dft_prbs_pass( dft_prbs_pass),
	.dll_core( dll_core),
	.dq_diff_in( dq_diff_in),
	.dq_sstl_in( dq_sstl_in),
	.dqs_diff_in_0( dqs_diff_in_0),
	.dqs_diff_in_1( dqs_diff_in_1),
	.dqs_diff_in_2( dqs_diff_in_2),
	.dqs_diff_in_3( dqs_diff_in_3),
	.dqs_sstl_n_0( dqs_sstl_n_0),
	.dqs_sstl_n_1( dqs_sstl_n_1),
	.dqs_sstl_n_2( dqs_sstl_n_2),
	.dqs_sstl_n_3( dqs_sstl_n_3),
	.dqs_sstl_p_0( dqs_sstl_p_0),
	.dqs_sstl_p_1( dqs_sstl_p_1),
	.dqs_sstl_p_2( dqs_sstl_p_2),
	.dqs_sstl_p_3( dqs_sstl_p_3),
	.dzoutx( dzoutx),
	.early_bhniotri( early_bhniotri),
	.early_csren( early_csren),
	.early_enrnsl( early_enrnsl),
	.early_frzreg( early_frzreg),
	.early_nfrzdrv( early_nfrzdrv),
	.early_niotri( early_niotri),
	.early_plniotri( early_plniotri),
	.early_usrmode( early_usrmode),
	.enrnsl( enrnsl),
	.entest( entest),
	.fb_clkout( fb_clkout),
	.fr_in_clk( fr_in_clk),
	.fr_out_clk( fr_out_clk),
	.frzreg( frzreg),
	.hps_to_core_ctrl_en( hps_to_core_ctrl_en),
	.hr_in_clk( hr_in_clk),
	.hr_out_clk( hr_out_clk),
	.i50u_ref( i50u_ref),
	.ibp50u( ibp50u),
	.ibp50u_cal( ibp50u_cal),
	.ioereg_locked( ioereg_locked),
	.jtag_clk( jtag_clk),
	.jtag_highz( jtag_highz),
	.jtag_mode( jtag_mode),
	.jtag_sdin( jtag_sdin),
	.jtag_sdout( jtag_sdout),
	.jtag_shftdr( jtag_shftdr),
	.jtag_updtdr( jtag_updtdr),
	.lane_cal_done( lane_cal_done),
	.local_bhniotri( local_bhniotri),
	.local_enrnsl( local_enrnsl),
	.local_frzreg( local_frzreg),
	.local_nfrzdrv( local_nfrzdrv),
	.local_niotri( local_niotri),
	.local_plniotri( local_plniotri),
	.local_usrmode( local_usrmode),
	.local_wkpullup( local_wkpullup),
	.lvds_rx_clk_chnl0( lvds_rx_clk_chnl0),
	.lvds_rx_clk_chnl1( lvds_rx_clk_chnl1),
	.lvds_rx_clk_chnl2( lvds_rx_clk_chnl2),
	.lvds_rx_clk_chnl3( lvds_rx_clk_chnl3),
	.lvds_rx_clk_chnl4( lvds_rx_clk_chnl4),
	.lvds_rx_clk_chnl5( lvds_rx_clk_chnl5),
	.lvds_tx_clk_chnl0( lvds_tx_clk_chnl0),
	.lvds_tx_clk_chnl1( lvds_tx_clk_chnl1),
	.lvds_tx_clk_chnl2( lvds_tx_clk_chnl2),
	.lvds_tx_clk_chnl3( lvds_tx_clk_chnl3),
	.lvds_tx_clk_chnl4( lvds_tx_clk_chnl4),
	.lvds_tx_clk_chnl5( lvds_tx_clk_chnl5),
	.mrnk_read_core( mrnk_read_core),
	.mrnk_write_core( mrnk_write_core),
	.n_crnt_clk( n_crnt_clk),
	.n_next_clk( n_next_clk),
	.naclr( naclr),
	.ncein( ncein),
	.nceout( nceout),
	.next_clk( next_clk),
	.nfrzdrv( nfrzdrv),
	.niotri( niotri),
	.nsclr( nsclr),
	.oct_enable( oct_enable),
	.oeb_from_core( oeb_from_core),
	.osc_en_n( osc_en_n),
	.osc_enable_in( osc_enable_in),
	.osc_mode_in( osc_mode_in),
	.osc_rocount_to_core( osc_rocount_to_core),
	.osc_sel_n( osc_sel_n),
	.phy_clk( phy_clk),
	.phy_clk_phs( phy_clk_phs),
	.pipeline_global_en_n( pipeline_global_en_n),
	.pll_clk( pll_clk),
	.pll_locked( pll_locked),
	.plniotri( plniotri),
	.progctl( progctl),
	.progoe( progoe),
	.progout( progout),
	.rdata_en_full_core( rdata_en_full_core),
	.rdata_valid_core( rdata_valid_core),
	.regulator_clk( regulator_clk),
	.reinit( reinit),
	.reset_n( reset_n),
	.scan_shift_n( scan_shift_n),
	.scanin( scanin),
	.scanout( scanout),
	.switch_dn( switch_dn),
	.switch_up( switch_up),
	.sync_clk_bot_in( sync_clk_bot_in),
	.sync_clk_bot_out( sync_clk_bot_out),
	.sync_clk_top_in( sync_clk_top_in),
	.sync_clk_top_out( sync_clk_top_out),
	.sync_data_bot_in( sync_data_bot_in),
	.sync_data_bot_out( sync_data_bot_out),
	.sync_data_top_in( sync_data_top_in),
	.sync_data_top_out( sync_data_top_out),
	.test_avl_clk_in_en_n( test_avl_clk_in_en_n),
	.test_clk( test_clk),
	.test_clk_ph_buf_en_n( test_clk_ph_buf_en_n),
	.test_clk_pll_en_n( test_clk_pll_en_n),
	.test_clr_n( test_clr_n),
	.test_datovr_en_n( test_datovr_en_n),
	.test_db_csr_in( test_db_csr_in),
	.test_dbg_in( test_dbg_in),
	.test_dbg_out( test_dbg_out),
	.test_dqs_csr_in( test_dqs_csr_in),
	.test_dqs_enable_en_n( test_dqs_enable_en_n),
	.test_fr_clk_en_n( test_fr_clk_en_n),
	.test_hr_clk_en_n( test_hr_clk_en_n),
	.test_int_clk_en_n( test_int_clk_en_n),
	.test_interp_clk_en_n( test_interp_clk_en_n),
	.test_ioereg2_csr_out( test_ioereg2_csr_out),
	.test_phy_clk_en_n( test_phy_clk_en_n),
	.test_phy_clk_lane_en_n( test_phy_clk_lane_en_n),
	.test_pst_clk_en_n( test_pst_clk_en_n),
	.test_pst_dll_i( test_pst_dll_i),
	.test_pst_dll_o( test_pst_dll_o),
	.test_tdf_select_n( test_tdf_select_n),
	.test_vref_csr_out( test_vref_csr_out),
	.test_xor_clk( test_xor_clk),
	.tpctl( tpctl),
	.tpdata( tpdata),
	.tpin( tpin),
	.up_ph( up_ph),
	.usrmode( usrmode),
	.vref_ext( vref_ext),
	.vref_int( vref_int),
	.weak_pullup_enable( weak_pullup_enable),
	.wkpullup( wkpullup),
	.x1024_osc_out( x1024_osc_out),
	.xor_vref( xor_vref),
	.xprio_clk( xprio_clk),
	.xprio_sync( xprio_sync),
	.xprio_xbus( xprio_xbus)
);

endmodule
