//
// Wrapper for CSR read and write structures and functions.
//

`ifndef CCI_CSR_IF_VH
`define CCI_CSR_IF_VH

import cci_csr_if_pkg::*;
import ccip_feature_list_pkg::*;

`endif
