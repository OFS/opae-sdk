// ed_sim_clks_sharing_splitter.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module ed_sim_clks_sharing_splitter (
		input  wire [31:0] sig_input,    //    sig_input_if.clks_sharing
		output wire [31:0] sig_output_0  // sig_output_if_0.clks_sharing
	);

	assign sig_output_0 = sig_input;

endmodule
