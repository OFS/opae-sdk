//
// Wrapper for MPF shim structures and functions.
//

`ifndef CCI_MPF_SHIM_VH
`define CCI_MPF_SHIM_VH

import cci_mpf_shim_pkg::*;

`endif
